module miniRISC (clk,
    sys_rst,
    din,
    dout);
 input clk;
 input sys_rst;
 input [15:0] din;
 output [15:0] dout;

 wire \GPR[0][0] ;
 wire \GPR[0][10] ;
 wire \GPR[0][11] ;
 wire \GPR[0][12] ;
 wire \GPR[0][13] ;
 wire \GPR[0][14] ;
 wire \GPR[0][15] ;
 wire \GPR[0][1] ;
 wire \GPR[0][2] ;
 wire \GPR[0][3] ;
 wire \GPR[0][4] ;
 wire \GPR[0][5] ;
 wire \GPR[0][6] ;
 wire \GPR[0][7] ;
 wire \GPR[0][8] ;
 wire \GPR[0][9] ;
 wire \GPR[1][0] ;
 wire \GPR[1][10] ;
 wire \GPR[1][11] ;
 wire \GPR[1][12] ;
 wire \GPR[1][13] ;
 wire \GPR[1][14] ;
 wire \GPR[1][15] ;
 wire \GPR[1][1] ;
 wire \GPR[1][2] ;
 wire \GPR[1][3] ;
 wire \GPR[1][4] ;
 wire \GPR[1][5] ;
 wire \GPR[1][6] ;
 wire \GPR[1][7] ;
 wire \GPR[1][8] ;
 wire \GPR[1][9] ;
 wire \GPR[2][0] ;
 wire \GPR[2][10] ;
 wire \GPR[2][11] ;
 wire \GPR[2][12] ;
 wire \GPR[2][13] ;
 wire \GPR[2][14] ;
 wire \GPR[2][15] ;
 wire \GPR[2][1] ;
 wire \GPR[2][2] ;
 wire \GPR[2][3] ;
 wire \GPR[2][4] ;
 wire \GPR[2][5] ;
 wire \GPR[2][6] ;
 wire \GPR[2][7] ;
 wire \GPR[2][8] ;
 wire \GPR[2][9] ;
 wire \GPR[3][0] ;
 wire \GPR[3][10] ;
 wire \GPR[3][11] ;
 wire \GPR[3][12] ;
 wire \GPR[3][13] ;
 wire \GPR[3][14] ;
 wire \GPR[3][15] ;
 wire \GPR[3][1] ;
 wire \GPR[3][2] ;
 wire \GPR[3][3] ;
 wire \GPR[3][4] ;
 wire \GPR[3][5] ;
 wire \GPR[3][6] ;
 wire \GPR[3][7] ;
 wire \GPR[3][8] ;
 wire \GPR[3][9] ;
 wire \IR[0] ;
 wire clknet_3_7__leaf_clk;
 wire \IR[16] ;
 wire \IR[17] ;
 wire \IR[18] ;
 wire \IR[1] ;
 wire \IR[22] ;
 wire \IR[23] ;
 wire \IR[24] ;
 wire \IR[27] ;
 wire \IR[28] ;
 wire \IR[2] ;
 wire \IR[30] ;
 wire net35;
 wire \PC[0] ;
 wire \PC[1] ;
 wire \PC[2] ;
 wire \PC[3] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0918_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire jmp_flag;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire stop;
 wire zero;
 wire net;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_0__leaf_clk;
 wire net48;
 wire net47;
 wire net42;
 wire clknet_0_clk;
 wire net49;
 wire net46;
 wire net45;
 wire net44;
 wire net43;

 sky130_fd_sc_hd__edfxtp_1 \GPR[0][0]$_DFFE_PP_  (.D(_0000_),
    .DE(net42),
    .Q(\GPR[0][0] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][10]$_DFFE_PP_  (.D(_0001_),
    .DE(_0016_),
    .Q(\GPR[0][10] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][11]$_DFFE_PP_  (.D(_0002_),
    .DE(_0016_),
    .Q(\GPR[0][11] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][12]$_DFFE_PP_  (.D(_0003_),
    .DE(_0016_),
    .Q(\GPR[0][12] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][13]$_DFFE_PP_  (.D(_0004_),
    .DE(_0016_),
    .Q(\GPR[0][13] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][14]$_DFFE_PP_  (.D(_0005_),
    .DE(_0016_),
    .Q(\GPR[0][14] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][15]$_DFFE_PP_  (.D(_0006_),
    .DE(_0016_),
    .Q(\GPR[0][15] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][1]$_DFFE_PP_  (.D(_0007_),
    .DE(net42),
    .Q(\GPR[0][1] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][2]$_DFFE_PP_  (.D(_0008_),
    .DE(net42),
    .Q(\GPR[0][2] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][3]$_DFFE_PP_  (.D(_0009_),
    .DE(net42),
    .Q(\GPR[0][3] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][4]$_DFFE_PP_  (.D(_0010_),
    .DE(net42),
    .Q(\GPR[0][4] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][5]$_DFFE_PP_  (.D(_0011_),
    .DE(net42),
    .Q(\GPR[0][5] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][6]$_DFFE_PP_  (.D(_0012_),
    .DE(net42),
    .Q(\GPR[0][6] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][7]$_DFFE_PP_  (.D(_0013_),
    .DE(net42),
    .Q(\GPR[0][7] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][8]$_DFFE_PP_  (.D(_0014_),
    .DE(net42),
    .Q(\GPR[0][8] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[0][9]$_DFFE_PP_  (.D(_0015_),
    .DE(net42),
    .Q(\GPR[0][9] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][0]$_DFFE_PP_  (.D(_0000_),
    .DE(net43),
    .Q(\GPR[1][0] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][10]$_DFFE_PP_  (.D(_0001_),
    .DE(net43),
    .Q(\GPR[1][10] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][11]$_DFFE_PP_  (.D(_0002_),
    .DE(net43),
    .Q(\GPR[1][11] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][12]$_DFFE_PP_  (.D(_0003_),
    .DE(net43),
    .Q(\GPR[1][12] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][13]$_DFFE_PP_  (.D(_0004_),
    .DE(net43),
    .Q(\GPR[1][13] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][14]$_DFFE_PP_  (.D(_0005_),
    .DE(net43),
    .Q(\GPR[1][14] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][15]$_DFFE_PP_  (.D(_0006_),
    .DE(net43),
    .Q(\GPR[1][15] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][1]$_DFFE_PP_  (.D(_0007_),
    .DE(net43),
    .Q(\GPR[1][1] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][2]$_DFFE_PP_  (.D(_0008_),
    .DE(net43),
    .Q(\GPR[1][2] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][3]$_DFFE_PP_  (.D(_0009_),
    .DE(net43),
    .Q(\GPR[1][3] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][4]$_DFFE_PP_  (.D(_0010_),
    .DE(net43),
    .Q(\GPR[1][4] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][5]$_DFFE_PP_  (.D(_0011_),
    .DE(net43),
    .Q(\GPR[1][5] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][6]$_DFFE_PP_  (.D(_0012_),
    .DE(net43),
    .Q(\GPR[1][6] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][7]$_DFFE_PP_  (.D(_0013_),
    .DE(net43),
    .Q(\GPR[1][7] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][8]$_DFFE_PP_  (.D(_0014_),
    .DE(net43),
    .Q(\GPR[1][8] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[1][9]$_DFFE_PP_  (.D(_0015_),
    .DE(net43),
    .Q(\GPR[1][9] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][0]$_DFFE_PP_  (.D(_0000_),
    .DE(_0018_),
    .Q(\GPR[2][0] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][10]$_DFFE_PP_  (.D(_0001_),
    .DE(_0018_),
    .Q(\GPR[2][10] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][11]$_DFFE_PP_  (.D(_0002_),
    .DE(_0018_),
    .Q(\GPR[2][11] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][12]$_DFFE_PP_  (.D(_0003_),
    .DE(_0018_),
    .Q(\GPR[2][12] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][13]$_DFFE_PP_  (.D(_0004_),
    .DE(_0018_),
    .Q(\GPR[2][13] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][14]$_DFFE_PP_  (.D(_0005_),
    .DE(_0018_),
    .Q(\GPR[2][14] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][15]$_DFFE_PP_  (.D(_0006_),
    .DE(_0018_),
    .Q(\GPR[2][15] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][1]$_DFFE_PP_  (.D(_0007_),
    .DE(net44),
    .Q(\GPR[2][1] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][2]$_DFFE_PP_  (.D(_0008_),
    .DE(net44),
    .Q(\GPR[2][2] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][3]$_DFFE_PP_  (.D(_0009_),
    .DE(net44),
    .Q(\GPR[2][3] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][4]$_DFFE_PP_  (.D(_0010_),
    .DE(net44),
    .Q(\GPR[2][4] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][5]$_DFFE_PP_  (.D(_0011_),
    .DE(net44),
    .Q(\GPR[2][5] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][6]$_DFFE_PP_  (.D(_0012_),
    .DE(net44),
    .Q(\GPR[2][6] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][7]$_DFFE_PP_  (.D(_0013_),
    .DE(net44),
    .Q(\GPR[2][7] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][8]$_DFFE_PP_  (.D(_0014_),
    .DE(net44),
    .Q(\GPR[2][8] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[2][9]$_DFFE_PP_  (.D(_0015_),
    .DE(net44),
    .Q(\GPR[2][9] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][0]$_DFFE_PP_  (.D(_0000_),
    .DE(net45),
    .Q(\GPR[3][0] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][10]$_DFFE_PP_  (.D(_0001_),
    .DE(net45),
    .Q(\GPR[3][10] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][11]$_DFFE_PP_  (.D(_0002_),
    .DE(net45),
    .Q(\GPR[3][11] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][12]$_DFFE_PP_  (.D(_0003_),
    .DE(net45),
    .Q(\GPR[3][12] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][13]$_DFFE_PP_  (.D(_0004_),
    .DE(net45),
    .Q(\GPR[3][13] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][14]$_DFFE_PP_  (.D(_0005_),
    .DE(net45),
    .Q(\GPR[3][14] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][15]$_DFFE_PP_  (.D(_0006_),
    .DE(net45),
    .Q(\GPR[3][15] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][1]$_DFFE_PP_  (.D(_0007_),
    .DE(net45),
    .Q(\GPR[3][1] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][2]$_DFFE_PP_  (.D(_0008_),
    .DE(net45),
    .Q(\GPR[3][2] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][3]$_DFFE_PP_  (.D(_0009_),
    .DE(net45),
    .Q(\GPR[3][3] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][4]$_DFFE_PP_  (.D(_0010_),
    .DE(net45),
    .Q(\GPR[3][4] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][5]$_DFFE_PP_  (.D(_0011_),
    .DE(net45),
    .Q(\GPR[3][5] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][6]$_DFFE_PP_  (.D(_0012_),
    .DE(net45),
    .Q(\GPR[3][6] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][7]$_DFFE_PP_  (.D(_0013_),
    .DE(net45),
    .Q(\GPR[3][7] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][8]$_DFFE_PP_  (.D(_0014_),
    .DE(net45),
    .Q(\GPR[3][8] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \GPR[3][9]$_DFFE_PP_  (.D(_0015_),
    .DE(net45),
    .Q(\GPR[3][9] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[0]$_SDFFE_PP0P_  (.D(_0146_),
    .Q(\IR[0] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[16]$_SDFFE_PP0P_  (.D(_0147_),
    .Q(\IR[16] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[17]$_SDFFE_PP0P_  (.D(_0148_),
    .Q(\IR[17] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[18]$_SDFFE_PP0P_  (.D(_0149_),
    .Q(\IR[18] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[1]$_SDFFE_PP0P_  (.D(_0150_),
    .Q(\IR[1] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[22]$_SDFFE_PP0P_  (.D(_0151_),
    .Q(\IR[22] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[23]$_SDFFE_PP0P_  (.D(_0152_),
    .Q(\IR[23] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[24]$_SDFFE_PP0P_  (.D(_0153_),
    .Q(\IR[24] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[27]$_SDFFE_PP0P_  (.D(_0154_),
    .Q(\IR[27] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[28]$_SDFFE_PP0P_  (.D(_0155_),
    .Q(\IR[28] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[2]$_SDFFE_PP0P_  (.D(_0156_),
    .Q(\IR[2] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \IR[30]$_SDFFE_PP0P_  (.D(_0157_),
    .Q(\IR[30] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \PC[0]$_SDFFE_PP0P_  (.D(_0158_),
    .Q(\PC[0] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \PC[1]$_SDFFE_PP0P_  (.D(_0159_),
    .Q(\PC[1] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \PC[2]$_SDFFE_PP0P_  (.D(_0160_),
    .Q(\PC[2] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \PC[3]$_SDFFE_PP0P_  (.D(_0161_),
    .Q(\PC[3] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__inv_1 _0959_ (.A(\IR[23] ),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_1 _0960_ (.A(\IR[27] ),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_1 _0961_ (.A(net35),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_1 _0962_ (.A(\IR[30] ),
    .Y(_0275_));
 sky130_fd_sc_hd__inv_1 _0964_ (.A(\state[1] ),
    .Y(_0277_));
 sky130_fd_sc_hd__nor3_2 _0965_ (.A(\state[2] ),
    .B(\state[0] ),
    .C(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__o2111ai_1 _0966_ (.A1(\IR[28] ),
    .A2(_0273_),
    .B1(_0274_),
    .C1(_0275_),
    .D1(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__nand2_1 _0967_ (.A(_0278_),
    .B(_0274_),
    .Y(_0280_));
 sky130_fd_sc_hd__nor2_1 _0968_ (.A(\IR[16] ),
    .B(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__nor3_1 _0969_ (.A(\IR[30] ),
    .B(\IR[28] ),
    .C(_0273_),
    .Y(_0282_));
 sky130_fd_sc_hd__nand2_1 _0970_ (.A(_0281_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_1 _0972_ (.A(\IR[16] ),
    .Y(_0285_));
 sky130_fd_sc_hd__nor2_1 _0973_ (.A(_0285_),
    .B(_0280_),
    .Y(_0286_));
 sky130_fd_sc_hd__nand2_1 _0974_ (.A(_0286_),
    .B(_0282_),
    .Y(_0287_));
 sky130_fd_sc_hd__nand3_1 _0975_ (.A(_0279_),
    .B(_0283_),
    .C(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__nand3b_1 _0976_ (.A_N(\IR[24] ),
    .B(_0288_),
    .C(\IR[22] ),
    .Y(_0289_));
 sky130_fd_sc_hd__nor2_2 _0977_ (.A(_0272_),
    .B(_0289_),
    .Y(_0019_));
 sky130_fd_sc_hd__nor2_1 _0978_ (.A(\IR[22] ),
    .B(\IR[24] ),
    .Y(_0290_));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(_0288_),
    .B(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__nor2_2 _0980_ (.A(_0272_),
    .B(_0291_),
    .Y(_0018_));
 sky130_fd_sc_hd__nor2_2 _0981_ (.A(\IR[23] ),
    .B(_0289_),
    .Y(_0017_));
 sky130_fd_sc_hd__nor2_2 _0982_ (.A(\IR[23] ),
    .B(_0291_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_1 _0985_ (.A(\GPR[0][14] ),
    .Y(_0129_));
 sky130_fd_sc_hd__a21oi_1 _0989_ (.A1(net49),
    .A2(\GPR[1][14] ),
    .B1(net48),
    .Y(_0297_));
 sky130_fd_sc_hd__o21ai_0 _0990_ (.A1(net49),
    .A2(_0129_),
    .B1(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__inv_2 _0991_ (.A(net49),
    .Y(_0299_));
 sky130_fd_sc_hd__nand2_1 _0993_ (.A(_0299_),
    .B(\GPR[2][14] ),
    .Y(_0301_));
 sky130_fd_sc_hd__nand2_1 _0994_ (.A(net49),
    .B(\GPR[3][14] ),
    .Y(_0302_));
 sky130_fd_sc_hd__nand3_1 _0995_ (.A(_0301_),
    .B(net48),
    .C(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__nand2_1 _0996_ (.A(_0298_),
    .B(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_1 _0997_ (.A(_0304_),
    .Y(_0128_));
 sky130_fd_sc_hd__nand2_1 _0998_ (.A(_0299_),
    .B(\GPR[2][13] ),
    .Y(_0305_));
 sky130_fd_sc_hd__nand2_1 _1000_ (.A(net49),
    .B(\GPR[3][13] ),
    .Y(_0307_));
 sky130_fd_sc_hd__nand3_1 _1001_ (.A(_0305_),
    .B(net48),
    .C(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__nand2_1 _1002_ (.A(_0299_),
    .B(\GPR[0][13] ),
    .Y(_0309_));
 sky130_fd_sc_hd__inv_2 _1003_ (.A(\IR[18] ),
    .Y(_0310_));
 sky130_fd_sc_hd__nand2_1 _1005_ (.A(net49),
    .B(\GPR[1][13] ),
    .Y(_0312_));
 sky130_fd_sc_hd__nand3_1 _1006_ (.A(_0309_),
    .B(_0310_),
    .C(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__nand2_1 _1007_ (.A(_0308_),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__inv_2 _1008_ (.A(_0314_),
    .Y(_0122_));
 sky130_fd_sc_hd__nand2_1 _1010_ (.A(_0299_),
    .B(\GPR[2][12] ),
    .Y(_0316_));
 sky130_fd_sc_hd__nand2_1 _1011_ (.A(net49),
    .B(\GPR[3][12] ),
    .Y(_0317_));
 sky130_fd_sc_hd__nand3_1 _1012_ (.A(_0316_),
    .B(net48),
    .C(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__nand2_1 _1013_ (.A(_0299_),
    .B(\GPR[0][12] ),
    .Y(_0319_));
 sky130_fd_sc_hd__nand2_1 _1014_ (.A(net49),
    .B(\GPR[1][12] ),
    .Y(_0320_));
 sky130_fd_sc_hd__nand3_1 _1015_ (.A(_0319_),
    .B(_0310_),
    .C(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__nand2_2 _1016_ (.A(_0318_),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_1 _1017_ (.A(_0322_),
    .Y(_0116_));
 sky130_fd_sc_hd__nand2_1 _1018_ (.A(_0299_),
    .B(\GPR[2][11] ),
    .Y(_0323_));
 sky130_fd_sc_hd__nand2_1 _1019_ (.A(net49),
    .B(\GPR[3][11] ),
    .Y(_0324_));
 sky130_fd_sc_hd__nand3_1 _1020_ (.A(_0323_),
    .B(net48),
    .C(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__nand2_1 _1021_ (.A(_0299_),
    .B(\GPR[0][11] ),
    .Y(_0326_));
 sky130_fd_sc_hd__nand2_1 _1022_ (.A(net49),
    .B(\GPR[1][11] ),
    .Y(_0327_));
 sky130_fd_sc_hd__nand3_1 _1023_ (.A(_0326_),
    .B(_0310_),
    .C(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__nand2_2 _1024_ (.A(_0325_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__inv_2 _1025_ (.A(_0329_),
    .Y(_0110_));
 sky130_fd_sc_hd__nand2_1 _1026_ (.A(_0299_),
    .B(\GPR[0][10] ),
    .Y(_0330_));
 sky130_fd_sc_hd__nand2_1 _1027_ (.A(net49),
    .B(\GPR[1][10] ),
    .Y(_0331_));
 sky130_fd_sc_hd__nand2_1 _1028_ (.A(_0330_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__nand2_1 _1030_ (.A(_0332_),
    .B(_0310_),
    .Y(_0334_));
 sky130_fd_sc_hd__nand2_1 _1031_ (.A(_0299_),
    .B(\GPR[2][10] ),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _1032_ (.A(net49),
    .B(\GPR[3][10] ),
    .Y(_0336_));
 sky130_fd_sc_hd__nand2_1 _1033_ (.A(_0335_),
    .B(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__nand2_1 _1034_ (.A(_0337_),
    .B(net48),
    .Y(_0338_));
 sky130_fd_sc_hd__nand2_1 _1035_ (.A(_0334_),
    .B(_0338_),
    .Y(_0104_));
 sky130_fd_sc_hd__nand2_1 _1037_ (.A(_0299_),
    .B(\GPR[0][9] ),
    .Y(_0340_));
 sky130_fd_sc_hd__nand2_1 _1038_ (.A(net49),
    .B(\GPR[1][9] ),
    .Y(_0341_));
 sky130_fd_sc_hd__nand2_1 _1039_ (.A(_0340_),
    .B(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_1 _1040_ (.A(_0342_),
    .B(_0310_),
    .Y(_0343_));
 sky130_fd_sc_hd__nand2_1 _1041_ (.A(_0299_),
    .B(\GPR[2][9] ),
    .Y(_0344_));
 sky130_fd_sc_hd__nand2_1 _1042_ (.A(net49),
    .B(\GPR[3][9] ),
    .Y(_0345_));
 sky130_fd_sc_hd__nand2_1 _1043_ (.A(_0344_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__nand2_1 _1044_ (.A(_0346_),
    .B(net48),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _1045_ (.A(_0343_),
    .B(_0347_),
    .Y(_0098_));
 sky130_fd_sc_hd__nand2_1 _1046_ (.A(_0299_),
    .B(\GPR[0][8] ),
    .Y(_0348_));
 sky130_fd_sc_hd__nand2_1 _1047_ (.A(net49),
    .B(\GPR[1][8] ),
    .Y(_0349_));
 sky130_fd_sc_hd__nand2_1 _1048_ (.A(_0348_),
    .B(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_1 _1049_ (.A(_0350_),
    .B(_0310_),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_1 _1050_ (.A(_0299_),
    .B(\GPR[2][8] ),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _1051_ (.A(net49),
    .B(\GPR[3][8] ),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_1 _1052_ (.A(_0352_),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__nand2_1 _1053_ (.A(_0354_),
    .B(net48),
    .Y(_0355_));
 sky130_fd_sc_hd__nand2_1 _1054_ (.A(_0351_),
    .B(_0355_),
    .Y(_0092_));
 sky130_fd_sc_hd__nand2_1 _1055_ (.A(_0299_),
    .B(\GPR[2][7] ),
    .Y(_0356_));
 sky130_fd_sc_hd__nand2_1 _1056_ (.A(net49),
    .B(\GPR[3][7] ),
    .Y(_0357_));
 sky130_fd_sc_hd__nand3_1 _1057_ (.A(_0356_),
    .B(net48),
    .C(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_1 _1058_ (.A(_0299_),
    .B(\GPR[0][7] ),
    .Y(_0359_));
 sky130_fd_sc_hd__nand2_1 _1059_ (.A(net49),
    .B(\GPR[1][7] ),
    .Y(_0360_));
 sky130_fd_sc_hd__nand3_2 _1060_ (.A(_0359_),
    .B(_0310_),
    .C(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2_2 _1061_ (.A(_0358_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(_0362_),
    .Y(_0086_));
 sky130_fd_sc_hd__nand2_1 _1063_ (.A(_0299_),
    .B(\GPR[2][6] ),
    .Y(_0363_));
 sky130_fd_sc_hd__nand2_1 _1064_ (.A(net49),
    .B(\GPR[3][6] ),
    .Y(_0364_));
 sky130_fd_sc_hd__nand3_1 _1065_ (.A(_0363_),
    .B(net48),
    .C(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__nand2_1 _1066_ (.A(_0299_),
    .B(\GPR[0][6] ),
    .Y(_0366_));
 sky130_fd_sc_hd__nand2_1 _1067_ (.A(net49),
    .B(\GPR[1][6] ),
    .Y(_0367_));
 sky130_fd_sc_hd__nand3_1 _1068_ (.A(_0366_),
    .B(_0310_),
    .C(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2_2 _1069_ (.A(_0365_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__inv_2 _1070_ (.A(_0369_),
    .Y(_0080_));
 sky130_fd_sc_hd__nand2_1 _1071_ (.A(_0299_),
    .B(\GPR[0][5] ),
    .Y(_0370_));
 sky130_fd_sc_hd__nand2_1 _1072_ (.A(net49),
    .B(\GPR[1][5] ),
    .Y(_0371_));
 sky130_fd_sc_hd__nand2_1 _1073_ (.A(_0370_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__nand2_1 _1074_ (.A(_0372_),
    .B(_0310_),
    .Y(_0373_));
 sky130_fd_sc_hd__nand2_1 _1075_ (.A(_0299_),
    .B(\GPR[2][5] ),
    .Y(_0374_));
 sky130_fd_sc_hd__nand2_1 _1076_ (.A(net49),
    .B(\GPR[3][5] ),
    .Y(_0375_));
 sky130_fd_sc_hd__nand2_1 _1077_ (.A(_0374_),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__nand2_1 _1078_ (.A(_0376_),
    .B(net48),
    .Y(_0377_));
 sky130_fd_sc_hd__nand2_1 _1079_ (.A(_0373_),
    .B(_0377_),
    .Y(_0074_));
 sky130_fd_sc_hd__nand2_1 _1080_ (.A(_0299_),
    .B(\GPR[0][4] ),
    .Y(_0378_));
 sky130_fd_sc_hd__nand2_1 _1081_ (.A(net49),
    .B(\GPR[1][4] ),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _1082_ (.A(_0378_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__nand2_1 _1083_ (.A(_0380_),
    .B(_0310_),
    .Y(_0381_));
 sky130_fd_sc_hd__inv_1 _1084_ (.A(\GPR[2][4] ),
    .Y(_0382_));
 sky130_fd_sc_hd__nand2_1 _1085_ (.A(_0299_),
    .B(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__inv_1 _1086_ (.A(\GPR[3][4] ),
    .Y(_0384_));
 sky130_fd_sc_hd__nand2_1 _1087_ (.A(_0384_),
    .B(net49),
    .Y(_0385_));
 sky130_fd_sc_hd__nand3_1 _1088_ (.A(_0383_),
    .B(_0385_),
    .C(net48),
    .Y(_0386_));
 sky130_fd_sc_hd__nand2_2 _1089_ (.A(_0381_),
    .B(_0386_),
    .Y(_0068_));
 sky130_fd_sc_hd__nand2_1 _1090_ (.A(_0299_),
    .B(\GPR[0][3] ),
    .Y(_0387_));
 sky130_fd_sc_hd__nand2_1 _1091_ (.A(net49),
    .B(\GPR[1][3] ),
    .Y(_0388_));
 sky130_fd_sc_hd__nand2_1 _1092_ (.A(_0387_),
    .B(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__nand2_1 _1093_ (.A(_0389_),
    .B(_0310_),
    .Y(_0390_));
 sky130_fd_sc_hd__inv_1 _1094_ (.A(\GPR[2][3] ),
    .Y(_0391_));
 sky130_fd_sc_hd__nand2_1 _1095_ (.A(_0299_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__inv_1 _1096_ (.A(\GPR[3][3] ),
    .Y(_0393_));
 sky130_fd_sc_hd__nand2_1 _1097_ (.A(_0393_),
    .B(net49),
    .Y(_0394_));
 sky130_fd_sc_hd__nand3_1 _1098_ (.A(_0392_),
    .B(_0394_),
    .C(net48),
    .Y(_0395_));
 sky130_fd_sc_hd__nand2_1 _1099_ (.A(_0390_),
    .B(_0395_),
    .Y(_0062_));
 sky130_fd_sc_hd__nor2_1 _1100_ (.A(\GPR[3][2] ),
    .B(_0299_),
    .Y(_0396_));
 sky130_fd_sc_hd__o21ai_0 _1101_ (.A1(net49),
    .A2(\GPR[2][2] ),
    .B1(net48),
    .Y(_0397_));
 sky130_fd_sc_hd__nor2_1 _1102_ (.A(net49),
    .B(\GPR[0][2] ),
    .Y(_0398_));
 sky130_fd_sc_hd__o21ai_0 _1103_ (.A1(\GPR[1][2] ),
    .A2(_0299_),
    .B1(_0310_),
    .Y(_0399_));
 sky130_fd_sc_hd__o22ai_1 _1104_ (.A1(_0396_),
    .A2(_0397_),
    .B1(_0398_),
    .B2(_0399_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_1 _1105_ (.A(\GPR[0][1] ),
    .Y(_0029_));
 sky130_fd_sc_hd__nor2_1 _1106_ (.A(net49),
    .B(_0029_),
    .Y(_0400_));
 sky130_fd_sc_hd__inv_1 _1107_ (.A(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__nand2_1 _1108_ (.A(net49),
    .B(\GPR[1][1] ),
    .Y(_0402_));
 sky130_fd_sc_hd__a21oi_1 _1109_ (.A1(net49),
    .A2(\GPR[3][1] ),
    .B1(_0310_),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _1110_ (.A(_0299_),
    .B(\GPR[2][1] ),
    .Y(_0404_));
 sky130_fd_sc_hd__a32oi_1 _1111_ (.A1(_0401_),
    .A2(_0402_),
    .A3(_0310_),
    .B1(_0403_),
    .B2(_0404_),
    .Y(_0020_));
 sky130_fd_sc_hd__nand2_1 _1112_ (.A(_0299_),
    .B(\GPR[0][0] ),
    .Y(_0405_));
 sky130_fd_sc_hd__nand2_1 _1113_ (.A(net49),
    .B(\GPR[1][0] ),
    .Y(_0406_));
 sky130_fd_sc_hd__a21oi_1 _1114_ (.A1(net49),
    .A2(\GPR[3][0] ),
    .B1(_0310_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand2_1 _1115_ (.A(_0299_),
    .B(\GPR[2][0] ),
    .Y(_0408_));
 sky130_fd_sc_hd__a32oi_1 _1116_ (.A1(_0405_),
    .A2(_0406_),
    .A3(_0310_),
    .B1(_0407_),
    .B2(_0408_),
    .Y(_0040_));
 sky130_fd_sc_hd__nand3_1 _1117_ (.A(_0275_),
    .B(\IR[27] ),
    .C(\IR[28] ),
    .Y(_0409_));
 sky130_fd_sc_hd__inv_1 _1118_ (.A(_0286_),
    .Y(_0410_));
 sky130_fd_sc_hd__nor2_1 _1119_ (.A(_0409_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__inv_2 _1120_ (.A(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__inv_1 _1122_ (.A(_0278_),
    .Y(_0414_));
 sky130_fd_sc_hd__nor4_1 _1123_ (.A(net35),
    .B(\IR[16] ),
    .C(_0409_),
    .D(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__inv_1 _1124_ (.A(net46),
    .Y(_0416_));
 sky130_fd_sc_hd__inv_1 _1125_ (.A(_0041_),
    .Y(_0417_));
 sky130_fd_sc_hd__nand2_1 _1126_ (.A(_0275_),
    .B(\IR[28] ),
    .Y(_0418_));
 sky130_fd_sc_hd__nor2_1 _1127_ (.A(\IR[27] ),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__inv_1 _1128_ (.A(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__inv_1 _1129_ (.A(_0281_),
    .Y(_0421_));
 sky130_fd_sc_hd__nor2_4 _1130_ (.A(_0420_),
    .B(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__nand2_1 _1131_ (.A(_0286_),
    .B(_0419_),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_1 _1132_ (.A(_0040_),
    .Y(_0038_));
 sky130_fd_sc_hd__nand3_1 _1133_ (.A(_0286_),
    .B(\IR[0] ),
    .C(_0282_),
    .Y(_0424_));
 sky130_fd_sc_hd__o221ai_1 _1134_ (.A1(_0039_),
    .A2(_0423_),
    .B1(_0283_),
    .B2(_0038_),
    .C1(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__a21oi_1 _1135_ (.A1(_0417_),
    .A2(_0422_),
    .B1(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__o221ai_1 _1136_ (.A1(_0042_),
    .A2(_0412_),
    .B1(_0043_),
    .B2(_0416_),
    .C1(_0426_),
    .Y(_0000_));
 sky130_fd_sc_hd__nor2_1 _1137_ (.A(_0409_),
    .B(_0421_),
    .Y(_0427_));
 sky130_fd_sc_hd__inv_1 _1138_ (.A(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_1 _1139_ (.A(\IR[1] ),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_1 _1140_ (.A(_0423_),
    .Y(_0429_));
 sky130_fd_sc_hd__nand2_1 _1141_ (.A(_0429_),
    .B(_0023_),
    .Y(_0430_));
 sky130_fd_sc_hd__nand2_1 _1142_ (.A(_0422_),
    .B(_0028_),
    .Y(_0431_));
 sky130_fd_sc_hd__inv_1 _1143_ (.A(_0283_),
    .Y(_0432_));
 sky130_fd_sc_hd__nand2_1 _1144_ (.A(net47),
    .B(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__o2111a_1 _1145_ (.A1(_0025_),
    .A2(_0287_),
    .B1(_0430_),
    .C1(_0431_),
    .D1(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__o221ai_1 _1146_ (.A1(_0032_),
    .A2(_0412_),
    .B1(_0035_),
    .B2(_0428_),
    .C1(_0434_),
    .Y(_0007_));
 sky130_fd_sc_hd__xnor2_1 _1147_ (.A(_0022_),
    .B(_0057_),
    .Y(_0435_));
 sky130_fd_sc_hd__inv_1 _1148_ (.A(\IR[2] ),
    .Y(_0055_));
 sky130_fd_sc_hd__nand2_1 _1149_ (.A(_0432_),
    .B(_0052_),
    .Y(_0436_));
 sky130_fd_sc_hd__o21ai_0 _1150_ (.A1(_0055_),
    .A2(_0287_),
    .B1(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__a21oi_1 _1151_ (.A1(_0429_),
    .A2(_0435_),
    .B1(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__xor2_1 _1152_ (.A(_0027_),
    .B(_0054_),
    .X(_0439_));
 sky130_fd_sc_hd__nand2_1 _1153_ (.A(_0422_),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__inv_1 _1154_ (.A(_0031_),
    .Y(_0441_));
 sky130_fd_sc_hd__nand2_1 _1155_ (.A(_0441_),
    .B(_0057_),
    .Y(_0442_));
 sky130_fd_sc_hd__inv_1 _1156_ (.A(_0057_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand2_1 _1157_ (.A(_0443_),
    .B(_0031_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand3_1 _1158_ (.A(_0411_),
    .B(_0442_),
    .C(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__xnor2_1 _1159_ (.A(_0034_),
    .B(_0061_),
    .Y(_0446_));
 sky130_fd_sc_hd__nand2_1 _1160_ (.A(net46),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__nand4_1 _1161_ (.A(_0438_),
    .B(_0440_),
    .C(_0445_),
    .D(_0447_),
    .Y(_0008_));
 sky130_fd_sc_hd__a21oi_1 _1162_ (.A1(_0050_),
    .A2(_0061_),
    .B1(_0060_),
    .Y(_0448_));
 sky130_fd_sc_hd__nand3b_1 _1163_ (.A_N(_0033_),
    .B(_0051_),
    .C(_0061_),
    .Y(_0449_));
 sky130_fd_sc_hd__nand2_1 _1164_ (.A(_0448_),
    .B(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__xnor2_1 _1165_ (.A(_0067_),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__nand2_1 _1166_ (.A(_0057_),
    .B(_0048_),
    .Y(_0452_));
 sky130_fd_sc_hd__inv_1 _1167_ (.A(_0056_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand2_1 _1168_ (.A(_0452_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__nand2_1 _1169_ (.A(_0057_),
    .B(_0049_),
    .Y(_0455_));
 sky130_fd_sc_hd__nor2_1 _1170_ (.A(_0030_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__o21ai_0 _1171_ (.A1(_0454_),
    .A2(_0456_),
    .B1(_0062_),
    .Y(_0457_));
 sky130_fd_sc_hd__nand2_1 _1172_ (.A(_0299_),
    .B(\GPR[2][3] ),
    .Y(_0458_));
 sky130_fd_sc_hd__nand2_1 _1173_ (.A(net49),
    .B(\GPR[3][3] ),
    .Y(_0459_));
 sky130_fd_sc_hd__nand3_2 _1174_ (.A(_0458_),
    .B(net48),
    .C(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__nand3_2 _1175_ (.A(_0387_),
    .B(_0310_),
    .C(_0388_),
    .Y(_0461_));
 sky130_fd_sc_hd__nand2_2 _1176_ (.A(_0460_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__nor2_1 _1177_ (.A(_0454_),
    .B(_0456_),
    .Y(_0463_));
 sky130_fd_sc_hd__nand2_1 _1178_ (.A(_0462_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__nand2_1 _1179_ (.A(_0457_),
    .B(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__clkinv_1 _1180_ (.A(_0422_),
    .Y(_0466_));
 sky130_fd_sc_hd__a21oi_1 _1181_ (.A1(_0046_),
    .A2(_0054_),
    .B1(_0053_),
    .Y(_0467_));
 sky130_fd_sc_hd__nand3_1 _1182_ (.A(_0026_),
    .B(_0047_),
    .C(_0054_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2_1 _1183_ (.A(_0467_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__xnor2_1 _1184_ (.A(_0064_),
    .B(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand3_1 _1185_ (.A(_0443_),
    .B(_0021_),
    .C(_0045_),
    .Y(_0471_));
 sky130_fd_sc_hd__inv_1 _1186_ (.A(_0058_),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2_1 _1187_ (.A(_0443_),
    .B(_0044_),
    .Y(_0473_));
 sky130_fd_sc_hd__nand3_1 _1188_ (.A(_0471_),
    .B(_0472_),
    .C(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2_1 _1189_ (.A(_0462_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__nand2_1 _1190_ (.A(_0473_),
    .B(_0472_),
    .Y(_0476_));
 sky130_fd_sc_hd__inv_1 _1191_ (.A(_0471_),
    .Y(_0477_));
 sky130_fd_sc_hd__nor2_1 _1192_ (.A(_0476_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__nand2_1 _1193_ (.A(_0062_),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__a21oi_1 _1194_ (.A1(_0475_),
    .A2(_0479_),
    .B1(_0423_),
    .Y(_0480_));
 sky130_fd_sc_hd__a21oi_1 _1195_ (.A1(_0432_),
    .A2(_0062_),
    .B1(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__o21ai_1 _1196_ (.A1(_0466_),
    .A2(_0470_),
    .B1(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__a21oi_1 _1197_ (.A1(_0411_),
    .A2(_0465_),
    .B1(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__o21ai_0 _1198_ (.A1(_0428_),
    .A2(_0451_),
    .B1(_0483_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_1 _1199_ (.A(_0073_),
    .Y(_0484_));
 sky130_fd_sc_hd__a21oi_1 _1200_ (.A1(_0060_),
    .A2(_0067_),
    .B1(_0066_),
    .Y(_0485_));
 sky130_fd_sc_hd__inv_1 _1201_ (.A(_0034_),
    .Y(_0486_));
 sky130_fd_sc_hd__nand3_1 _1202_ (.A(_0486_),
    .B(_0061_),
    .C(_0067_),
    .Y(_0487_));
 sky130_fd_sc_hd__nand2_1 _1203_ (.A(_0485_),
    .B(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__xor2_1 _1204_ (.A(_0484_),
    .B(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nand2_1 _1205_ (.A(_0299_),
    .B(\GPR[2][4] ),
    .Y(_0490_));
 sky130_fd_sc_hd__nand2_1 _1206_ (.A(net49),
    .B(\GPR[3][4] ),
    .Y(_0491_));
 sky130_fd_sc_hd__nand3_1 _1207_ (.A(_0490_),
    .B(net48),
    .C(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__nand3_1 _1208_ (.A(_0378_),
    .B(_0310_),
    .C(_0379_),
    .Y(_0493_));
 sky130_fd_sc_hd__nand2_4 _1209_ (.A(_0492_),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__nand2_1 _1210_ (.A(_0443_),
    .B(_0022_),
    .Y(_0495_));
 sky130_fd_sc_hd__nand2_1 _1211_ (.A(_0495_),
    .B(_0472_),
    .Y(_0496_));
 sky130_fd_sc_hd__nand3_1 _1212_ (.A(_0062_),
    .B(_0494_),
    .C(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__nand3_1 _1213_ (.A(_0460_),
    .B(_0461_),
    .C(_0496_),
    .Y(_0498_));
 sky130_fd_sc_hd__nand2_1 _1214_ (.A(_0498_),
    .B(_0068_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _1215_ (.A(_0497_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__nor2_1 _1216_ (.A(_0494_),
    .B(_0283_),
    .Y(_0501_));
 sky130_fd_sc_hd__inv_1 _1217_ (.A(_0070_),
    .Y(_0502_));
 sky130_fd_sc_hd__a21oi_1 _1218_ (.A1(_0053_),
    .A2(_0064_),
    .B1(_0063_),
    .Y(_0503_));
 sky130_fd_sc_hd__nand3_1 _1219_ (.A(_0027_),
    .B(_0054_),
    .C(_0064_),
    .Y(_0504_));
 sky130_fd_sc_hd__nand2_1 _1220_ (.A(_0503_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__xor2_1 _1221_ (.A(_0502_),
    .B(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__nor2_1 _1222_ (.A(_0506_),
    .B(_0466_),
    .Y(_0507_));
 sky130_fd_sc_hd__nand3_1 _1223_ (.A(_0462_),
    .B(_0453_),
    .C(_0442_),
    .Y(_0508_));
 sky130_fd_sc_hd__inv_2 _1224_ (.A(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__nand2_1 _1225_ (.A(_0509_),
    .B(_0068_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand2_1 _1226_ (.A(_0508_),
    .B(_0494_),
    .Y(_0511_));
 sky130_fd_sc_hd__nand2_1 _1227_ (.A(_0510_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__nor2_1 _1228_ (.A(_0412_),
    .B(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__a2111oi_0 _1229_ (.A1(_0429_),
    .A2(_0500_),
    .B1(_0501_),
    .C1(_0507_),
    .D1(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__o21ai_0 _1230_ (.A1(_0416_),
    .A2(_0489_),
    .B1(_0514_),
    .Y(_0010_));
 sky130_fd_sc_hd__nand2_1 _1231_ (.A(_0064_),
    .B(_0070_),
    .Y(_0515_));
 sky130_fd_sc_hd__inv_1 _1232_ (.A(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__nand2_1 _1233_ (.A(_0469_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__nand2_1 _1234_ (.A(_0063_),
    .B(_0070_),
    .Y(_0518_));
 sky130_fd_sc_hd__inv_1 _1235_ (.A(_0069_),
    .Y(_0519_));
 sky130_fd_sc_hd__nand2_1 _1236_ (.A(_0518_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__inv_1 _1237_ (.A(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _1238_ (.A(_0517_),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__xor2_1 _1239_ (.A(_0076_),
    .B(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__nand3_1 _1240_ (.A(_0374_),
    .B(net48),
    .C(_0375_),
    .Y(_0524_));
 sky130_fd_sc_hd__nand3_2 _1241_ (.A(_0370_),
    .B(_0310_),
    .C(_0371_),
    .Y(_0525_));
 sky130_fd_sc_hd__nand2_4 _1242_ (.A(_0524_),
    .B(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__nor2_2 _1243_ (.A(_0478_),
    .B(_0462_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand2_1 _1244_ (.A(_0527_),
    .B(_0068_),
    .Y(_0528_));
 sky130_fd_sc_hd__nand2_1 _1245_ (.A(_0528_),
    .B(_0526_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand3_1 _1246_ (.A(_0527_),
    .B(_0074_),
    .C(_0068_),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _1247_ (.A(_0529_),
    .B(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__o22ai_1 _1248_ (.A1(_0283_),
    .A2(_0526_),
    .B1(_0423_),
    .B2(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__a21oi_1 _1249_ (.A1(_0422_),
    .A2(_0523_),
    .B1(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__nand3_2 _1250_ (.A(_0494_),
    .B(_0462_),
    .C(_0463_),
    .Y(_0534_));
 sky130_fd_sc_hd__xor2_1 _1251_ (.A(_0526_),
    .B(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__nand2_1 _1252_ (.A(_0535_),
    .B(_0411_),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_1 _1253_ (.A(_0067_),
    .B(_0073_),
    .Y(_0537_));
 sky130_fd_sc_hd__inv_1 _1254_ (.A(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__nand2_1 _1255_ (.A(_0450_),
    .B(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _1256_ (.A(_0066_),
    .B(_0073_),
    .Y(_0540_));
 sky130_fd_sc_hd__inv_1 _1257_ (.A(_0072_),
    .Y(_0541_));
 sky130_fd_sc_hd__nand2_1 _1258_ (.A(_0540_),
    .B(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__inv_1 _1259_ (.A(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__nand2_1 _1260_ (.A(_0539_),
    .B(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__xor2_1 _1261_ (.A(_0079_),
    .B(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__nand2_1 _1262_ (.A(_0545_),
    .B(_0427_),
    .Y(_0546_));
 sky130_fd_sc_hd__nand3_1 _1263_ (.A(_0533_),
    .B(_0536_),
    .C(_0546_),
    .Y(_0011_));
 sky130_fd_sc_hd__nand2_2 _1264_ (.A(_0526_),
    .B(_0494_),
    .Y(_0547_));
 sky130_fd_sc_hd__o21ai_0 _1265_ (.A1(_0547_),
    .A2(_0508_),
    .B1(_0369_),
    .Y(_0548_));
 sky130_fd_sc_hd__nor2_1 _1266_ (.A(_0547_),
    .B(_0508_),
    .Y(_0549_));
 sky130_fd_sc_hd__nand2_1 _1267_ (.A(_0549_),
    .B(_0080_),
    .Y(_0550_));
 sky130_fd_sc_hd__nand2_1 _1268_ (.A(_0548_),
    .B(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__nand2_1 _1269_ (.A(_0061_),
    .B(_0067_),
    .Y(_0552_));
 sky130_fd_sc_hd__nand2_1 _1270_ (.A(_0073_),
    .B(_0079_),
    .Y(_0553_));
 sky130_fd_sc_hd__nor3_1 _1271_ (.A(_0034_),
    .B(_0552_),
    .C(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__a21oi_1 _1272_ (.A1(_0072_),
    .A2(_0079_),
    .B1(_0078_),
    .Y(_0555_));
 sky130_fd_sc_hd__o21ai_0 _1273_ (.A1(_0553_),
    .A2(_0485_),
    .B1(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__nor2_1 _1274_ (.A(_0554_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__xor2_1 _1275_ (.A(_0085_),
    .B(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__nand2_1 _1276_ (.A(_0070_),
    .B(_0076_),
    .Y(_0559_));
 sky130_fd_sc_hd__inv_1 _1277_ (.A(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__nand2_1 _1278_ (.A(_0505_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__a21oi_1 _1279_ (.A1(_0069_),
    .A2(_0076_),
    .B1(_0075_),
    .Y(_0562_));
 sky130_fd_sc_hd__nand2_1 _1280_ (.A(_0561_),
    .B(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__xor2_1 _1281_ (.A(_0082_),
    .B(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__nand2_1 _1282_ (.A(_0074_),
    .B(_0068_),
    .Y(_0565_));
 sky130_fd_sc_hd__nor2_1 _1283_ (.A(_0498_),
    .B(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__nand2_1 _1284_ (.A(_0566_),
    .B(_0369_),
    .Y(_0567_));
 sky130_fd_sc_hd__nor2_8 _1285_ (.A(_0526_),
    .B(_0494_),
    .Y(_0568_));
 sky130_fd_sc_hd__inv_1 _1286_ (.A(_0498_),
    .Y(_0569_));
 sky130_fd_sc_hd__nand2_2 _1287_ (.A(_0568_),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_1 _1288_ (.A(_0570_),
    .B(_0080_),
    .Y(_0571_));
 sky130_fd_sc_hd__nand2_1 _1289_ (.A(_0567_),
    .B(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__nor2_1 _1290_ (.A(_0369_),
    .B(_0283_),
    .Y(_0573_));
 sky130_fd_sc_hd__a221oi_1 _1291_ (.A1(_0564_),
    .A2(_0422_),
    .B1(_0572_),
    .B2(_0429_),
    .C1(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__o221ai_1 _1292_ (.A1(_0412_),
    .A2(_0551_),
    .B1(_0428_),
    .B2(_0558_),
    .C1(_0574_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_1 _1293_ (.A(_0091_),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2_1 _1294_ (.A(_0079_),
    .B(_0085_),
    .Y(_0576_));
 sky130_fd_sc_hd__inv_1 _1295_ (.A(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__nand3_1 _1296_ (.A(_0450_),
    .B(_0538_),
    .C(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__a21oi_1 _1297_ (.A1(_0078_),
    .A2(_0085_),
    .B1(_0084_),
    .Y(_0579_));
 sky130_fd_sc_hd__inv_1 _1298_ (.A(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__a21oi_1 _1299_ (.A1(_0542_),
    .A2(_0577_),
    .B1(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_1 _1300_ (.A(_0578_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__xor2_1 _1301_ (.A(_0575_),
    .B(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__nand2_1 _1302_ (.A(_0076_),
    .B(_0082_),
    .Y(_0584_));
 sky130_fd_sc_hd__inv_1 _1303_ (.A(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__nand3_1 _1304_ (.A(_0469_),
    .B(_0516_),
    .C(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__nand2_1 _1305_ (.A(_0075_),
    .B(_0082_),
    .Y(_0587_));
 sky130_fd_sc_hd__inv_1 _1306_ (.A(_0081_),
    .Y(_0588_));
 sky130_fd_sc_hd__nand2_1 _1307_ (.A(_0587_),
    .B(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__a21oi_1 _1308_ (.A1(_0520_),
    .A2(_0585_),
    .B1(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _1309_ (.A(_0586_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__xor2_1 _1310_ (.A(_0088_),
    .B(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__nand2_2 _1311_ (.A(_0369_),
    .B(_0526_),
    .Y(_0593_));
 sky130_fd_sc_hd__o21ai_0 _1312_ (.A1(_0593_),
    .A2(_0534_),
    .B1(_0362_),
    .Y(_0594_));
 sky130_fd_sc_hd__nor2_1 _1313_ (.A(_0593_),
    .B(_0534_),
    .Y(_0595_));
 sky130_fd_sc_hd__nand2_1 _1314_ (.A(_0595_),
    .B(_0086_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _1315_ (.A(_0594_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__nor2_1 _1316_ (.A(_0412_),
    .B(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__nand3_2 _1317_ (.A(_0568_),
    .B(_0527_),
    .C(_0080_),
    .Y(_0599_));
 sky130_fd_sc_hd__nand2_1 _1318_ (.A(_0599_),
    .B(_0086_),
    .Y(_0600_));
 sky130_fd_sc_hd__nand3_1 _1319_ (.A(_0474_),
    .B(_0460_),
    .C(_0461_),
    .Y(_0601_));
 sky130_fd_sc_hd__nor2_1 _1320_ (.A(_0369_),
    .B(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand3_1 _1321_ (.A(_0602_),
    .B(_0362_),
    .C(_0568_),
    .Y(_0603_));
 sky130_fd_sc_hd__nand2_1 _1322_ (.A(_0600_),
    .B(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__nand2_1 _1323_ (.A(_0604_),
    .B(_0429_),
    .Y(_0605_));
 sky130_fd_sc_hd__o21ai_0 _1324_ (.A1(_0283_),
    .A2(_0362_),
    .B1(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__a211oi_1 _1325_ (.A1(_0422_),
    .A2(_0592_),
    .B1(_0598_),
    .C1(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__o21ai_0 _1326_ (.A1(_0416_),
    .A2(_0583_),
    .B1(_0607_),
    .Y(_0013_));
 sky130_fd_sc_hd__nand2_1 _1327_ (.A(_0362_),
    .B(_0369_),
    .Y(_0608_));
 sky130_fd_sc_hd__nor2_2 _1328_ (.A(_0547_),
    .B(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__nand2_1 _1329_ (.A(_0609_),
    .B(_0509_),
    .Y(_0610_));
 sky130_fd_sc_hd__nand3_1 _1330_ (.A(_0352_),
    .B(net48),
    .C(_0353_),
    .Y(_0611_));
 sky130_fd_sc_hd__nand3_2 _1331_ (.A(_0348_),
    .B(_0310_),
    .C(_0349_),
    .Y(_0612_));
 sky130_fd_sc_hd__nand2_2 _1332_ (.A(_0611_),
    .B(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__nand2_1 _1333_ (.A(_0610_),
    .B(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__nand3_1 _1334_ (.A(_0609_),
    .B(_0509_),
    .C(_0092_),
    .Y(_0615_));
 sky130_fd_sc_hd__nand2_1 _1335_ (.A(_0614_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__a21o_1 _1336_ (.A1(_0084_),
    .A2(_0091_),
    .B1(_0090_),
    .X(_0617_));
 sky130_fd_sc_hd__nand2_1 _1337_ (.A(_0085_),
    .B(_0091_),
    .Y(_0618_));
 sky130_fd_sc_hd__nor2_1 _1338_ (.A(_0618_),
    .B(_0555_),
    .Y(_0619_));
 sky130_fd_sc_hd__nor2_1 _1339_ (.A(_0617_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__nor2_1 _1340_ (.A(_0553_),
    .B(_0618_),
    .Y(_0621_));
 sky130_fd_sc_hd__nand2_1 _1341_ (.A(_0488_),
    .B(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__nand2_1 _1342_ (.A(_0620_),
    .B(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__xnor2_1 _1343_ (.A(_0097_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nor2_2 _1344_ (.A(_0362_),
    .B(_0369_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand3_1 _1345_ (.A(_0568_),
    .B(_0625_),
    .C(_0569_),
    .Y(_0626_));
 sky130_fd_sc_hd__nand2_1 _1346_ (.A(_0626_),
    .B(_0092_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand3_1 _1347_ (.A(_0566_),
    .B(_0613_),
    .C(_0625_),
    .Y(_0628_));
 sky130_fd_sc_hd__nand2_1 _1348_ (.A(_0627_),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__nand2_1 _1349_ (.A(_0081_),
    .B(_0088_),
    .Y(_0630_));
 sky130_fd_sc_hd__inv_1 _1350_ (.A(_0087_),
    .Y(_0631_));
 sky130_fd_sc_hd__nand2_1 _1351_ (.A(_0630_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__nand2_1 _1352_ (.A(_0082_),
    .B(_0088_),
    .Y(_0633_));
 sky130_fd_sc_hd__nor2_1 _1353_ (.A(_0633_),
    .B(_0562_),
    .Y(_0634_));
 sky130_fd_sc_hd__nor2_1 _1354_ (.A(_0632_),
    .B(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__nor2_1 _1355_ (.A(_0559_),
    .B(_0633_),
    .Y(_0636_));
 sky130_fd_sc_hd__nand2_1 _1356_ (.A(_0505_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__nand2_1 _1357_ (.A(_0635_),
    .B(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__xnor2_1 _1358_ (.A(_0094_),
    .B(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__nor2_1 _1359_ (.A(_0466_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__a221oi_1 _1360_ (.A1(_0432_),
    .A2(_0092_),
    .B1(_0629_),
    .B2(_0429_),
    .C1(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__o221ai_1 _1361_ (.A1(_0412_),
    .A2(_0616_),
    .B1(_0428_),
    .B2(_0624_),
    .C1(_0641_),
    .Y(_0014_));
 sky130_fd_sc_hd__nand2_1 _1362_ (.A(_0088_),
    .B(_0094_),
    .Y(_0642_));
 sky130_fd_sc_hd__nor2_1 _1363_ (.A(_0584_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__nand2_1 _1364_ (.A(_0522_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand3_1 _1365_ (.A(_0589_),
    .B(_0088_),
    .C(_0094_),
    .Y(_0645_));
 sky130_fd_sc_hd__a21oi_1 _1366_ (.A1(_0087_),
    .A2(_0094_),
    .B1(_0093_),
    .Y(_0646_));
 sky130_fd_sc_hd__nand3_1 _1367_ (.A(_0644_),
    .B(_0645_),
    .C(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2_1 _1368_ (.A(_0647_),
    .B(_0100_),
    .Y(_0648_));
 sky130_fd_sc_hd__inv_1 _1369_ (.A(_0100_),
    .Y(_0649_));
 sky130_fd_sc_hd__nand4_1 _1370_ (.A(_0644_),
    .B(_0649_),
    .C(_0645_),
    .D(_0646_),
    .Y(_0650_));
 sky130_fd_sc_hd__nand2_1 _1371_ (.A(_0648_),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__nor2_1 _1372_ (.A(_0466_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__nand2_1 _1373_ (.A(_0613_),
    .B(_0362_),
    .Y(_0653_));
 sky130_fd_sc_hd__nor2_4 _1374_ (.A(_0593_),
    .B(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__inv_2 _1375_ (.A(_0534_),
    .Y(_0655_));
 sky130_fd_sc_hd__nand2_1 _1376_ (.A(_0654_),
    .B(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__nand3_1 _1377_ (.A(_0344_),
    .B(net48),
    .C(_0345_),
    .Y(_0657_));
 sky130_fd_sc_hd__nand3_1 _1378_ (.A(_0340_),
    .B(_0310_),
    .C(_0341_),
    .Y(_0658_));
 sky130_fd_sc_hd__nand2_1 _1379_ (.A(_0657_),
    .B(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__nand2_1 _1380_ (.A(_0656_),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__nand3_1 _1381_ (.A(_0654_),
    .B(_0655_),
    .C(_0098_),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2_1 _1382_ (.A(_0660_),
    .B(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__nor2_1 _1383_ (.A(_0412_),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__nand2_1 _1384_ (.A(_0527_),
    .B(_0080_),
    .Y(_0664_));
 sky130_fd_sc_hd__nor2_2 _1385_ (.A(_0565_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__nor2_2 _1386_ (.A(_0613_),
    .B(_0362_),
    .Y(_0666_));
 sky130_fd_sc_hd__nand2_1 _1387_ (.A(_0665_),
    .B(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__nand2_1 _1388_ (.A(_0667_),
    .B(_0659_),
    .Y(_0668_));
 sky130_fd_sc_hd__nand3_1 _1389_ (.A(_0665_),
    .B(_0098_),
    .C(_0666_),
    .Y(_0669_));
 sky130_fd_sc_hd__nand2_1 _1390_ (.A(_0668_),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__o22ai_1 _1391_ (.A1(_0283_),
    .A2(_0659_),
    .B1(_0423_),
    .B2(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__nor3_1 _1392_ (.A(_0652_),
    .B(_0663_),
    .C(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__nand2_1 _1393_ (.A(_0091_),
    .B(_0097_),
    .Y(_0673_));
 sky130_fd_sc_hd__nor2_1 _1394_ (.A(_0576_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__a21oi_1 _1395_ (.A1(_0090_),
    .A2(_0097_),
    .B1(_0096_),
    .Y(_0675_));
 sky130_fd_sc_hd__o21ai_0 _1396_ (.A1(_0673_),
    .A2(_0579_),
    .B1(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__a21oi_1 _1397_ (.A1(_0544_),
    .A2(_0674_),
    .B1(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__inv_1 _1398_ (.A(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__inv_1 _1399_ (.A(_0103_),
    .Y(_0679_));
 sky130_fd_sc_hd__nand2_1 _1400_ (.A(_0678_),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__nand2_1 _1401_ (.A(_0677_),
    .B(_0103_),
    .Y(_0681_));
 sky130_fd_sc_hd__nand2_1 _1402_ (.A(_0680_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2_1 _1403_ (.A(_0682_),
    .B(_0427_),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _1404_ (.A(_0672_),
    .B(_0683_),
    .Y(_0015_));
 sky130_fd_sc_hd__nand2_1 _1405_ (.A(_0094_),
    .B(_0100_),
    .Y(_0684_));
 sky130_fd_sc_hd__nor2_1 _1406_ (.A(_0633_),
    .B(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__nand2_1 _1407_ (.A(_0563_),
    .B(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__inv_1 _1408_ (.A(_0684_),
    .Y(_0687_));
 sky130_fd_sc_hd__a21oi_1 _1409_ (.A1(_0093_),
    .A2(_0100_),
    .B1(_0099_),
    .Y(_0688_));
 sky130_fd_sc_hd__a21boi_0 _1410_ (.A1(_0632_),
    .A2(_0687_),
    .B1_N(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__nand2_1 _1411_ (.A(_0686_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__xnor2_1 _1412_ (.A(_0106_),
    .B(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__nor2_1 _1413_ (.A(_0466_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__nand3_1 _1414_ (.A(_0335_),
    .B(net48),
    .C(_0336_),
    .Y(_0693_));
 sky130_fd_sc_hd__nand3_2 _1415_ (.A(_0330_),
    .B(_0310_),
    .C(_0331_),
    .Y(_0694_));
 sky130_fd_sc_hd__nand2_1 _1416_ (.A(_0693_),
    .B(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__nand2_1 _1417_ (.A(_0098_),
    .B(_0092_),
    .Y(_0696_));
 sky130_fd_sc_hd__inv_2 _1418_ (.A(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__nand2_1 _1419_ (.A(_0697_),
    .B(_0625_),
    .Y(_0698_));
 sky130_fd_sc_hd__o21ai_0 _1420_ (.A1(_0570_),
    .A2(_0698_),
    .B1(_0695_),
    .Y(_0699_));
 sky130_fd_sc_hd__nor2_2 _1421_ (.A(_0570_),
    .B(_0698_),
    .Y(_0700_));
 sky130_fd_sc_hd__nand2_1 _1422_ (.A(_0700_),
    .B(_0104_),
    .Y(_0701_));
 sky130_fd_sc_hd__nand2_1 _1423_ (.A(_0699_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__o22ai_1 _1424_ (.A1(_0283_),
    .A2(_0695_),
    .B1(_0423_),
    .B2(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__nor2_1 _1425_ (.A(_0692_),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__inv_1 _1426_ (.A(_0547_),
    .Y(_0705_));
 sky130_fd_sc_hd__nor2_1 _1427_ (.A(_0442_),
    .B(_0062_),
    .Y(_0706_));
 sky130_fd_sc_hd__nand2_1 _1428_ (.A(_0705_),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__nand2_1 _1429_ (.A(_0659_),
    .B(_0613_),
    .Y(_0708_));
 sky130_fd_sc_hd__nor2_2 _1430_ (.A(_0608_),
    .B(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__nand2_1 _1431_ (.A(_0462_),
    .B(_0453_),
    .Y(_0710_));
 sky130_fd_sc_hd__nor2_1 _1432_ (.A(_0710_),
    .B(_0547_),
    .Y(_0711_));
 sky130_fd_sc_hd__nand4_1 _1433_ (.A(_0707_),
    .B(_0709_),
    .C(_0711_),
    .D(_0104_),
    .Y(_0712_));
 sky130_fd_sc_hd__nand3_1 _1434_ (.A(_0707_),
    .B(_0709_),
    .C(_0711_),
    .Y(_0713_));
 sky130_fd_sc_hd__nand2_1 _1435_ (.A(_0713_),
    .B(_0695_),
    .Y(_0714_));
 sky130_fd_sc_hd__nand3_1 _1436_ (.A(_0712_),
    .B(_0714_),
    .C(_0411_),
    .Y(_0715_));
 sky130_fd_sc_hd__nand2_1 _1437_ (.A(_0097_),
    .B(_0103_),
    .Y(_0716_));
 sky130_fd_sc_hd__nor2_1 _1438_ (.A(_0618_),
    .B(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__nand2_1 _1439_ (.A(_0556_),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__inv_1 _1440_ (.A(_0716_),
    .Y(_0719_));
 sky130_fd_sc_hd__a21o_1 _1441_ (.A1(_0096_),
    .A2(_0103_),
    .B1(_0102_),
    .X(_0720_));
 sky130_fd_sc_hd__a21oi_1 _1442_ (.A1(_0617_),
    .A2(_0719_),
    .B1(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__nor2_1 _1443_ (.A(_0552_),
    .B(_0553_),
    .Y(_0722_));
 sky130_fd_sc_hd__nand3_1 _1444_ (.A(_0722_),
    .B(_0717_),
    .C(_0486_),
    .Y(_0723_));
 sky130_fd_sc_hd__nand3_1 _1445_ (.A(_0718_),
    .B(_0721_),
    .C(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__xor2_1 _1446_ (.A(_0109_),
    .B(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__nand2_1 _1447_ (.A(_0725_),
    .B(_0427_),
    .Y(_0726_));
 sky130_fd_sc_hd__nand3_1 _1448_ (.A(_0704_),
    .B(_0715_),
    .C(_0726_),
    .Y(_0001_));
 sky130_fd_sc_hd__nand2_1 _1449_ (.A(_0100_),
    .B(_0106_),
    .Y(_0727_));
 sky130_fd_sc_hd__nor2_1 _1450_ (.A(_0642_),
    .B(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__nand2_1 _1451_ (.A(_0591_),
    .B(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__a21oi_1 _1452_ (.A1(_0099_),
    .A2(_0106_),
    .B1(_0105_),
    .Y(_0730_));
 sky130_fd_sc_hd__o21ai_0 _1453_ (.A1(_0727_),
    .A2(_0646_),
    .B1(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__inv_1 _1454_ (.A(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__nand3b_1 _1455_ (.A_N(_0112_),
    .B(_0729_),
    .C(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__nand2_1 _1456_ (.A(_0729_),
    .B(_0732_),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_1 _1457_ (.A(_0734_),
    .B(_0112_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_1 _1458_ (.A(_0695_),
    .B(_0659_),
    .Y(_0736_));
 sky130_fd_sc_hd__nand2_1 _1459_ (.A(_0666_),
    .B(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__o21ai_0 _1460_ (.A1(_0737_),
    .A2(_0599_),
    .B1(_0329_),
    .Y(_0738_));
 sky130_fd_sc_hd__nor2_2 _1461_ (.A(_0737_),
    .B(_0599_),
    .Y(_0739_));
 sky130_fd_sc_hd__nand2_1 _1462_ (.A(_0739_),
    .B(_0110_),
    .Y(_0740_));
 sky130_fd_sc_hd__nand2_1 _1463_ (.A(_0738_),
    .B(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__o22ai_1 _1464_ (.A1(_0283_),
    .A2(_0329_),
    .B1(_0423_),
    .B2(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__a31oi_1 _1465_ (.A1(_0422_),
    .A2(_0733_),
    .A3(_0735_),
    .B1(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__nand2_1 _1466_ (.A(_0695_),
    .B(_0659_),
    .Y(_0744_));
 sky130_fd_sc_hd__inv_1 _1467_ (.A(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__nand3_1 _1468_ (.A(_0654_),
    .B(_0655_),
    .C(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__nand2_1 _1469_ (.A(_0746_),
    .B(_0329_),
    .Y(_0747_));
 sky130_fd_sc_hd__nand4_1 _1470_ (.A(_0654_),
    .B(_0655_),
    .C(_0110_),
    .D(_0745_),
    .Y(_0748_));
 sky130_fd_sc_hd__nand3_1 _1471_ (.A(_0747_),
    .B(_0748_),
    .C(_0411_),
    .Y(_0749_));
 sky130_fd_sc_hd__nand2_1 _1472_ (.A(_0103_),
    .B(_0109_),
    .Y(_0750_));
 sky130_fd_sc_hd__nor2_1 _1473_ (.A(_0673_),
    .B(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__nand2_1 _1474_ (.A(_0582_),
    .B(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__a21oi_1 _1475_ (.A1(_0102_),
    .A2(_0109_),
    .B1(_0108_),
    .Y(_0753_));
 sky130_fd_sc_hd__o21ai_0 _1476_ (.A1(_0750_),
    .A2(_0675_),
    .B1(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__inv_1 _1477_ (.A(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__nand2_1 _1478_ (.A(_0752_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__xor2_1 _1479_ (.A(_0115_),
    .B(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__nand2_1 _1480_ (.A(_0757_),
    .B(_0427_),
    .Y(_0758_));
 sky130_fd_sc_hd__nand3_1 _1481_ (.A(_0743_),
    .B(_0749_),
    .C(_0758_),
    .Y(_0002_));
 sky130_fd_sc_hd__nand2_1 _1482_ (.A(_0106_),
    .B(_0112_),
    .Y(_0759_));
 sky130_fd_sc_hd__nor2_1 _1483_ (.A(_0684_),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__nand2_1 _1484_ (.A(_0105_),
    .B(_0112_),
    .Y(_0761_));
 sky130_fd_sc_hd__inv_1 _1485_ (.A(_0111_),
    .Y(_0762_));
 sky130_fd_sc_hd__nand2_1 _1486_ (.A(_0761_),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__o21bai_1 _1487_ (.A1(_0759_),
    .A2(_0688_),
    .B1_N(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__a21oi_1 _1488_ (.A1(_0638_),
    .A2(_0760_),
    .B1(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__xor2_1 _1489_ (.A(_0118_),
    .B(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__nor2_1 _1490_ (.A(_0466_),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__nand2_1 _1491_ (.A(_0329_),
    .B(_0695_),
    .Y(_0768_));
 sky130_fd_sc_hd__nor2_1 _1492_ (.A(_0708_),
    .B(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__nand3_1 _1493_ (.A(_0609_),
    .B(_0769_),
    .C(_0509_),
    .Y(_0770_));
 sky130_fd_sc_hd__nand2_1 _1494_ (.A(_0770_),
    .B(_0322_),
    .Y(_0771_));
 sky130_fd_sc_hd__nand4_1 _1495_ (.A(_0609_),
    .B(_0769_),
    .C(_0116_),
    .D(_0509_),
    .Y(_0772_));
 sky130_fd_sc_hd__nand2_1 _1496_ (.A(_0771_),
    .B(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__nor2_1 _1497_ (.A(_0412_),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__nand2_1 _1498_ (.A(_0086_),
    .B(_0080_),
    .Y(_0775_));
 sky130_fd_sc_hd__nor2_1 _1499_ (.A(_0565_),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__nand2_1 _1500_ (.A(_0110_),
    .B(_0104_),
    .Y(_0777_));
 sky130_fd_sc_hd__nor2_1 _1501_ (.A(_0696_),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__nand3_1 _1502_ (.A(_0776_),
    .B(_0778_),
    .C(_0569_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand2_1 _1503_ (.A(_0779_),
    .B(_0322_),
    .Y(_0780_));
 sky130_fd_sc_hd__nand4_1 _1504_ (.A(_0776_),
    .B(_0778_),
    .C(_0116_),
    .D(_0569_),
    .Y(_0781_));
 sky130_fd_sc_hd__nand2_1 _1505_ (.A(_0780_),
    .B(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__o22ai_1 _1506_ (.A1(_0283_),
    .A2(_0322_),
    .B1(_0423_),
    .B2(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__nor3_1 _1507_ (.A(_0767_),
    .B(_0774_),
    .C(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__nand2_1 _1508_ (.A(_0109_),
    .B(_0115_),
    .Y(_0785_));
 sky130_fd_sc_hd__nor2_1 _1509_ (.A(_0716_),
    .B(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__nand2_1 _1510_ (.A(_0623_),
    .B(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__a21o_1 _1511_ (.A1(_0108_),
    .A2(_0115_),
    .B1(_0114_),
    .X(_0788_));
 sky130_fd_sc_hd__a31oi_1 _1512_ (.A1(_0720_),
    .A2(_0109_),
    .A3(_0115_),
    .B1(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__nand2_1 _1513_ (.A(_0787_),
    .B(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__xor2_1 _1514_ (.A(_0121_),
    .B(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__nand2_1 _1515_ (.A(_0791_),
    .B(_0427_),
    .Y(_0792_));
 sky130_fd_sc_hd__nand2_1 _1516_ (.A(_0784_),
    .B(_0792_),
    .Y(_0003_));
 sky130_fd_sc_hd__nand2_1 _1517_ (.A(_0322_),
    .B(_0329_),
    .Y(_0793_));
 sky130_fd_sc_hd__nor2_1 _1518_ (.A(_0744_),
    .B(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__nand4_1 _1519_ (.A(_0654_),
    .B(_0794_),
    .C(_0655_),
    .D(_0122_),
    .Y(_0795_));
 sky130_fd_sc_hd__nand3_1 _1520_ (.A(_0654_),
    .B(_0794_),
    .C(_0655_),
    .Y(_0796_));
 sky130_fd_sc_hd__nand2_1 _1521_ (.A(_0796_),
    .B(_0314_),
    .Y(_0797_));
 sky130_fd_sc_hd__nand2_1 _1522_ (.A(_0795_),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__nand2_1 _1523_ (.A(_0115_),
    .B(_0121_),
    .Y(_0799_));
 sky130_fd_sc_hd__nor2_1 _1524_ (.A(_0750_),
    .B(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__a21oi_1 _1525_ (.A1(_0114_),
    .A2(_0121_),
    .B1(_0120_),
    .Y(_0801_));
 sky130_fd_sc_hd__o21ai_0 _1526_ (.A1(_0799_),
    .A2(_0753_),
    .B1(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__a21oi_1 _1527_ (.A1(_0676_),
    .A2(_0800_),
    .B1(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__nand3_1 _1528_ (.A(_0544_),
    .B(_0674_),
    .C(_0800_),
    .Y(_0804_));
 sky130_fd_sc_hd__nand2_1 _1529_ (.A(_0803_),
    .B(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__xor2_1 _1530_ (.A(_0127_),
    .B(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__nand2_1 _1531_ (.A(_0806_),
    .B(_0427_),
    .Y(_0807_));
 sky130_fd_sc_hd__inv_1 _1532_ (.A(_0124_),
    .Y(_0808_));
 sky130_fd_sc_hd__nand2_1 _1533_ (.A(_0112_),
    .B(_0118_),
    .Y(_0809_));
 sky130_fd_sc_hd__nor2_1 _1534_ (.A(_0727_),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__nand3_1 _1535_ (.A(_0522_),
    .B(_0643_),
    .C(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_1 _1536_ (.A(_0645_),
    .B(_0646_),
    .Y(_0812_));
 sky130_fd_sc_hd__a21oi_1 _1537_ (.A1(_0111_),
    .A2(_0118_),
    .B1(_0117_),
    .Y(_0813_));
 sky130_fd_sc_hd__o21ai_0 _1538_ (.A1(_0809_),
    .A2(_0730_),
    .B1(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__a21oi_1 _1539_ (.A1(_0812_),
    .A2(_0810_),
    .B1(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__nand2_1 _1540_ (.A(_0811_),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__xor2_1 _1541_ (.A(_0808_),
    .B(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__nor2_1 _1542_ (.A(_0466_),
    .B(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__nor2_2 _1543_ (.A(_0322_),
    .B(_0329_),
    .Y(_0819_));
 sky130_fd_sc_hd__nand2_1 _1544_ (.A(_0739_),
    .B(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__nand2_1 _1545_ (.A(_0820_),
    .B(_0314_),
    .Y(_0821_));
 sky130_fd_sc_hd__nand3_1 _1546_ (.A(_0739_),
    .B(_0122_),
    .C(_0819_),
    .Y(_0822_));
 sky130_fd_sc_hd__nand2_1 _1547_ (.A(_0821_),
    .B(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__o22ai_1 _1548_ (.A1(_0283_),
    .A2(_0314_),
    .B1(_0423_),
    .B2(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__nor2_1 _1549_ (.A(_0818_),
    .B(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__o211ai_1 _1550_ (.A1(_0412_),
    .A2(_0798_),
    .B1(_0807_),
    .C1(_0825_),
    .Y(_0004_));
 sky130_fd_sc_hd__nand2_1 _1551_ (.A(_0121_),
    .B(_0127_),
    .Y(_0826_));
 sky130_fd_sc_hd__nor2_1 _1552_ (.A(_0785_),
    .B(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__inv_1 _1553_ (.A(_0127_),
    .Y(_0828_));
 sky130_fd_sc_hd__a21oi_1 _1554_ (.A1(_0788_),
    .A2(_0121_),
    .B1(_0120_),
    .Y(_0829_));
 sky130_fd_sc_hd__o21bai_1 _1555_ (.A1(_0828_),
    .A2(_0829_),
    .B1_N(_0126_),
    .Y(_0830_));
 sky130_fd_sc_hd__a21oi_1 _1556_ (.A1(_0724_),
    .A2(_0827_),
    .B1(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__xor2_1 _1557_ (.A(_0132_),
    .B(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__a21oi_1 _1558_ (.A1(_0763_),
    .A2(_0118_),
    .B1(_0117_),
    .Y(_0833_));
 sky130_fd_sc_hd__o21bai_1 _1559_ (.A1(_0808_),
    .A2(_0833_),
    .B1_N(_0123_),
    .Y(_0834_));
 sky130_fd_sc_hd__inv_1 _1560_ (.A(_0118_),
    .Y(_0835_));
 sky130_fd_sc_hd__nor3_1 _1561_ (.A(_0835_),
    .B(_0808_),
    .C(_0759_),
    .Y(_0836_));
 sky130_fd_sc_hd__inv_1 _1562_ (.A(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__nor2_1 _1563_ (.A(_0837_),
    .B(_0689_),
    .Y(_0838_));
 sky130_fd_sc_hd__nor2_1 _1564_ (.A(_0834_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__nand3_1 _1565_ (.A(_0563_),
    .B(_0685_),
    .C(_0836_),
    .Y(_0840_));
 sky130_fd_sc_hd__nand2_1 _1566_ (.A(_0839_),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__inv_1 _1567_ (.A(_0131_),
    .Y(_0842_));
 sky130_fd_sc_hd__nand2_1 _1568_ (.A(_0841_),
    .B(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__nand3_1 _1569_ (.A(_0839_),
    .B(_0840_),
    .C(_0131_),
    .Y(_0844_));
 sky130_fd_sc_hd__nand2_1 _1570_ (.A(_0843_),
    .B(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__nor2_1 _1571_ (.A(_0466_),
    .B(_0845_),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_1 _1572_ (.A(_0314_),
    .B(_0322_),
    .Y(_0847_));
 sky130_fd_sc_hd__nor2_1 _1573_ (.A(_0768_),
    .B(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__nand4_1 _1574_ (.A(_0549_),
    .B(_0709_),
    .C(_0848_),
    .D(_0304_),
    .Y(_0849_));
 sky130_fd_sc_hd__nand3_1 _1575_ (.A(_0549_),
    .B(_0709_),
    .C(_0848_),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_1 _1576_ (.A(_0850_),
    .B(_0128_),
    .Y(_0851_));
 sky130_fd_sc_hd__a21oi_1 _1577_ (.A1(_0849_),
    .A2(_0851_),
    .B1(_0412_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand2_1 _1578_ (.A(_0819_),
    .B(_0122_),
    .Y(_0853_));
 sky130_fd_sc_hd__nor2_1 _1579_ (.A(_0695_),
    .B(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__nand2_1 _1580_ (.A(_0700_),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__nand2_1 _1581_ (.A(_0855_),
    .B(_0304_),
    .Y(_0856_));
 sky130_fd_sc_hd__nand3_1 _1582_ (.A(_0700_),
    .B(_0854_),
    .C(_0128_),
    .Y(_0857_));
 sky130_fd_sc_hd__nand2_1 _1583_ (.A(_0856_),
    .B(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__o22ai_1 _1584_ (.A1(_0283_),
    .A2(_0304_),
    .B1(_0423_),
    .B2(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__nor3_1 _1585_ (.A(_0846_),
    .B(_0852_),
    .C(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__o21ai_0 _1586_ (.A1(_0428_),
    .A2(_0832_),
    .B1(_0860_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_1 _1587_ (.A(\GPR[0][15] ),
    .Y(_0861_));
 sky130_fd_sc_hd__a21oi_1 _1588_ (.A1(\GPR[1][15] ),
    .A2(net49),
    .B1(net48),
    .Y(_0862_));
 sky130_fd_sc_hd__o21ai_1 _1589_ (.A1(_0861_),
    .A2(net49),
    .B1(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__nand2_1 _1590_ (.A(_0299_),
    .B(\GPR[2][15] ),
    .Y(_0864_));
 sky130_fd_sc_hd__nand2_1 _1591_ (.A(net49),
    .B(\GPR[3][15] ),
    .Y(_0865_));
 sky130_fd_sc_hd__nand3_1 _1592_ (.A(_0864_),
    .B(net48),
    .C(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__nand2_1 _1593_ (.A(_0863_),
    .B(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__inv_1 _1594_ (.A(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__nor2_1 _1595_ (.A(_0304_),
    .B(_0853_),
    .Y(_0869_));
 sky130_fd_sc_hd__inv_1 _1596_ (.A(_0737_),
    .Y(_0870_));
 sky130_fd_sc_hd__nand3_1 _1597_ (.A(_0869_),
    .B(_0665_),
    .C(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__nand2_1 _1598_ (.A(_0871_),
    .B(_0868_),
    .Y(_0872_));
 sky130_fd_sc_hd__nand4_1 _1599_ (.A(_0869_),
    .B(_0665_),
    .C(_0870_),
    .D(_0867_),
    .Y(_0873_));
 sky130_fd_sc_hd__nand2_1 _1600_ (.A(_0872_),
    .B(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__nand2_1 _1601_ (.A(_0842_),
    .B(_0124_),
    .Y(_0875_));
 sky130_fd_sc_hd__nor2_1 _1602_ (.A(_0809_),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__nand3_1 _1603_ (.A(_0591_),
    .B(_0728_),
    .C(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__a21oi_1 _1604_ (.A1(_0842_),
    .A2(_0123_),
    .B1(_0133_),
    .Y(_0878_));
 sky130_fd_sc_hd__o21ai_0 _1605_ (.A1(_0875_),
    .A2(_0813_),
    .B1(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__a21oi_1 _1606_ (.A1(_0731_),
    .A2(_0876_),
    .B1(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2_1 _1607_ (.A(_0877_),
    .B(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__xor2_1 _1608_ (.A(\GPR[0][15] ),
    .B(_0867_),
    .X(_0882_));
 sky130_fd_sc_hd__inv_1 _1609_ (.A(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__nand2_1 _1610_ (.A(_0881_),
    .B(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__nand3_1 _1611_ (.A(_0882_),
    .B(_0877_),
    .C(_0880_),
    .Y(_0885_));
 sky130_fd_sc_hd__nand2_1 _1612_ (.A(_0884_),
    .B(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__nor2_1 _1613_ (.A(_0466_),
    .B(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__a221oi_1 _1614_ (.A1(_0432_),
    .A2(_0868_),
    .B1(_0874_),
    .B2(_0429_),
    .C1(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__nand2_1 _1615_ (.A(_0304_),
    .B(_0314_),
    .Y(_0889_));
 sky130_fd_sc_hd__nor2_1 _1616_ (.A(_0793_),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__nor2_1 _1617_ (.A(_0653_),
    .B(_0744_),
    .Y(_0891_));
 sky130_fd_sc_hd__nand3_1 _1618_ (.A(_0595_),
    .B(_0890_),
    .C(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__nand2_1 _1619_ (.A(_0892_),
    .B(_0868_),
    .Y(_0893_));
 sky130_fd_sc_hd__nand4_1 _1620_ (.A(_0595_),
    .B(_0890_),
    .C(_0891_),
    .D(_0867_),
    .Y(_0894_));
 sky130_fd_sc_hd__nand2_1 _1621_ (.A(_0893_),
    .B(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__nand2_1 _1622_ (.A(_0895_),
    .B(_0411_),
    .Y(_0896_));
 sky130_fd_sc_hd__inv_1 _1623_ (.A(_0132_),
    .Y(_0897_));
 sky130_fd_sc_hd__nor3_1 _1624_ (.A(_0828_),
    .B(_0897_),
    .C(_0799_),
    .Y(_0898_));
 sky130_fd_sc_hd__nand2_1 _1625_ (.A(_0756_),
    .B(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_1 _1626_ (.A(_0126_),
    .B(_0132_),
    .Y(_0900_));
 sky130_fd_sc_hd__nor3_1 _1627_ (.A(_0828_),
    .B(_0897_),
    .C(_0801_),
    .Y(_0901_));
 sky130_fd_sc_hd__nor2_1 _1628_ (.A(_0130_),
    .B(_0901_),
    .Y(_0902_));
 sky130_fd_sc_hd__nand3_1 _1629_ (.A(_0899_),
    .B(_0900_),
    .C(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__nand2_1 _1630_ (.A(_0903_),
    .B(_0882_),
    .Y(_0904_));
 sky130_fd_sc_hd__nand4_1 _1631_ (.A(_0899_),
    .B(_0883_),
    .C(_0900_),
    .D(_0902_),
    .Y(_0905_));
 sky130_fd_sc_hd__nand3_1 _1632_ (.A(_0904_),
    .B(_0905_),
    .C(net46),
    .Y(_0906_));
 sky130_fd_sc_hd__nand3_1 _1633_ (.A(_0888_),
    .B(_0896_),
    .C(_0906_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_1 _1634_ (.A(net47),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_1 _1635_ (.A(\GPR[0][2] ),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_1 _1636_ (.A(\GPR[0][3] ),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_1 _1637_ (.A(\GPR[0][4] ),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_1 _1638_ (.A(\GPR[0][5] ),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_1 _1639_ (.A(\GPR[0][6] ),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_1 _1640_ (.A(\GPR[0][8] ),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_1 _1641_ (.A(\GPR[0][9] ),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_1 _1642_ (.A(\GPR[0][10] ),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_1 _1643_ (.A(\GPR[0][12] ),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_1 _1644_ (.A(\GPR[0][13] ),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_1 _1645_ (.A(\PC[0] ),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_1 _1646_ (.A(\PC[1] ),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_1 _1647_ (.A(\GPR[0][7] ),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_1 _1648_ (.A(\GPR[0][11] ),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_1 _1649_ (.A(_0140_),
    .Y(_0907_));
 sky130_fd_sc_hd__nand2_1 _1650_ (.A(_0277_),
    .B(\state[0] ),
    .Y(_0908_));
 sky130_fd_sc_hd__nor2_1 _1651_ (.A(\state[2] ),
    .B(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__inv_1 _1652_ (.A(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__nor2_1 _1653_ (.A(\PC[3] ),
    .B(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__inv_1 _1654_ (.A(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__a21oi_1 _1655_ (.A1(\PC[2] ),
    .A2(_0907_),
    .B1(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__o21ai_0 _1656_ (.A1(\PC[2] ),
    .A2(_0136_),
    .B1(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__nor2_1 _1657_ (.A(\state[2] ),
    .B(\state[1] ),
    .Y(_0915_));
 sky130_fd_sc_hd__inv_1 _1658_ (.A(_0915_),
    .Y(_0916_));
 sky130_fd_sc_hd__nand2_1 _1660_ (.A(_0916_),
    .B(\IR[0] ),
    .Y(_0918_));
 sky130_fd_sc_hd__a21oi_1 _1662_ (.A1(_0914_),
    .A2(_0918_),
    .B1(net35),
    .Y(_0146_));
 sky130_fd_sc_hd__a21oi_1 _1663_ (.A1(\IR[16] ),
    .A2(_0916_),
    .B1(_0913_),
    .Y(_0920_));
 sky130_fd_sc_hd__nor2_1 _1664_ (.A(net35),
    .B(_0920_),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_1 _1665_ (.A(\PC[2] ),
    .Y(_0921_));
 sky130_fd_sc_hd__nor2_1 _1666_ (.A(\PC[3] ),
    .B(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__inv_1 _1667_ (.A(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__nor3_1 _1668_ (.A(_0907_),
    .B(_0923_),
    .C(_0910_),
    .Y(_0924_));
 sky130_fd_sc_hd__a21oi_1 _1669_ (.A1(net49),
    .A2(_0916_),
    .B1(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__nor2_1 _1670_ (.A(net35),
    .B(_0925_),
    .Y(_0148_));
 sky130_fd_sc_hd__nor2_1 _1671_ (.A(_0139_),
    .B(_0923_),
    .Y(_0926_));
 sky130_fd_sc_hd__nand2_1 _1672_ (.A(_0926_),
    .B(_0909_),
    .Y(_0927_));
 sky130_fd_sc_hd__nand2_1 _1673_ (.A(_0916_),
    .B(net48),
    .Y(_0928_));
 sky130_fd_sc_hd__a21oi_1 _1674_ (.A1(_0927_),
    .A2(_0928_),
    .B1(net35),
    .Y(_0149_));
 sky130_fd_sc_hd__nor3_1 _1675_ (.A(_0134_),
    .B(\PC[2] ),
    .C(_0912_),
    .Y(_0929_));
 sky130_fd_sc_hd__a21oi_1 _1676_ (.A1(\IR[1] ),
    .A2(_0916_),
    .B1(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__nor2_1 _1677_ (.A(net35),
    .B(_0930_),
    .Y(_0150_));
 sky130_fd_sc_hd__nor2_1 _1678_ (.A(_0924_),
    .B(_0929_),
    .Y(_0931_));
 sky130_fd_sc_hd__nand2_1 _1679_ (.A(_0916_),
    .B(\IR[22] ),
    .Y(_0932_));
 sky130_fd_sc_hd__a21oi_1 _1680_ (.A1(_0931_),
    .A2(_0932_),
    .B1(net35),
    .Y(_0151_));
 sky130_fd_sc_hd__o22ai_1 _1681_ (.A1(_0272_),
    .A2(_0915_),
    .B1(_0144_),
    .B2(_0912_),
    .Y(_0933_));
 sky130_fd_sc_hd__inv_1 _1682_ (.A(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__nor2_1 _1683_ (.A(net35),
    .B(_0934_),
    .Y(_0152_));
 sky130_fd_sc_hd__nand2_1 _1684_ (.A(_0911_),
    .B(_0141_),
    .Y(_0935_));
 sky130_fd_sc_hd__nand2_1 _1685_ (.A(_0916_),
    .B(\IR[24] ),
    .Y(_0936_));
 sky130_fd_sc_hd__a21oi_1 _1686_ (.A1(_0935_),
    .A2(_0936_),
    .B1(net35),
    .Y(_0153_));
 sky130_fd_sc_hd__o21ai_0 _1687_ (.A1(\PC[0] ),
    .A2(_0923_),
    .B1(_0909_),
    .Y(_0937_));
 sky130_fd_sc_hd__nand2_1 _1688_ (.A(_0916_),
    .B(\IR[27] ),
    .Y(_0938_));
 sky130_fd_sc_hd__a21oi_1 _1689_ (.A1(_0937_),
    .A2(_0938_),
    .B1(net35),
    .Y(_0154_));
 sky130_fd_sc_hd__o21ai_0 _1690_ (.A1(\PC[3] ),
    .A2(_0143_),
    .B1(_0909_),
    .Y(_0939_));
 sky130_fd_sc_hd__nand2_1 _1691_ (.A(_0916_),
    .B(\IR[28] ),
    .Y(_0940_));
 sky130_fd_sc_hd__a21oi_1 _1692_ (.A1(_0939_),
    .A2(_0940_),
    .B1(net35),
    .Y(_0155_));
 sky130_fd_sc_hd__nand2_1 _1693_ (.A(\PC[2] ),
    .B(_0138_),
    .Y(_0941_));
 sky130_fd_sc_hd__o21ai_0 _1694_ (.A1(\PC[2] ),
    .A2(_0139_),
    .B1(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__a22oi_1 _1695_ (.A1(\IR[2] ),
    .A2(_0916_),
    .B1(_0911_),
    .B2(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__nor2_1 _1696_ (.A(net35),
    .B(_0943_),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_1 _1697_ (.A(\PC[3] ),
    .Y(_0944_));
 sky130_fd_sc_hd__nand2_1 _1698_ (.A(_0941_),
    .B(_0944_),
    .Y(_0171_));
 sky130_fd_sc_hd__nand2_1 _1699_ (.A(_0909_),
    .B(_0171_),
    .Y(_0172_));
 sky130_fd_sc_hd__nand2_1 _1700_ (.A(_0916_),
    .B(\IR[30] ),
    .Y(_0173_));
 sky130_fd_sc_hd__a21oi_1 _1701_ (.A1(_0172_),
    .A2(_0173_),
    .B1(net35),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_1 _1702_ (.A(\state[0] ),
    .Y(_0174_));
 sky130_fd_sc_hd__nor3_1 _1703_ (.A(\state[2] ),
    .B(_0174_),
    .C(_0277_),
    .Y(_0175_));
 sky130_fd_sc_hd__o21bai_1 _1704_ (.A1(\state[0] ),
    .A2(_0916_),
    .B1_N(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_1 _1705_ (.A(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__nand2_1 _1706_ (.A(_0177_),
    .B(\PC[0] ),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_1 _1707_ (.A(jmp_flag),
    .Y(_0179_));
 sky130_fd_sc_hd__nand2_1 _1708_ (.A(_0179_),
    .B(\PC[0] ),
    .Y(_0180_));
 sky130_fd_sc_hd__o211ai_1 _1709_ (.A1(\IR[0] ),
    .A2(_0179_),
    .B1(_0180_),
    .C1(_0175_),
    .Y(_0181_));
 sky130_fd_sc_hd__a21oi_1 _1710_ (.A1(_0178_),
    .A2(_0181_),
    .B1(net35),
    .Y(_0158_));
 sky130_fd_sc_hd__nand2_1 _1711_ (.A(_0177_),
    .B(\PC[1] ),
    .Y(_0182_));
 sky130_fd_sc_hd__nand2_1 _1712_ (.A(_0025_),
    .B(jmp_flag),
    .Y(_0183_));
 sky130_fd_sc_hd__o211ai_1 _1713_ (.A1(jmp_flag),
    .A2(_0137_),
    .B1(_0183_),
    .C1(_0175_),
    .Y(_0184_));
 sky130_fd_sc_hd__a21oi_1 _1714_ (.A1(_0182_),
    .A2(_0184_),
    .B1(net35),
    .Y(_0159_));
 sky130_fd_sc_hd__nand2_1 _1715_ (.A(_0177_),
    .B(\PC[2] ),
    .Y(_0185_));
 sky130_fd_sc_hd__nand2_1 _1716_ (.A(_0055_),
    .B(jmp_flag),
    .Y(_0186_));
 sky130_fd_sc_hd__o211ai_1 _1717_ (.A1(jmp_flag),
    .A2(_0142_),
    .B1(_0186_),
    .C1(_0175_),
    .Y(_0187_));
 sky130_fd_sc_hd__a21oi_1 _1718_ (.A1(_0185_),
    .A2(_0187_),
    .B1(net35),
    .Y(_0160_));
 sky130_fd_sc_hd__nand2_1 _1719_ (.A(_0177_),
    .B(\PC[3] ),
    .Y(_0188_));
 sky130_fd_sc_hd__nand2_1 _1720_ (.A(\PC[0] ),
    .B(_0145_),
    .Y(_0189_));
 sky130_fd_sc_hd__xor2_1 _1721_ (.A(_0944_),
    .B(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__nand3_1 _1722_ (.A(_0190_),
    .B(_0179_),
    .C(_0175_),
    .Y(_0191_));
 sky130_fd_sc_hd__a21oi_1 _1723_ (.A1(_0188_),
    .A2(_0191_),
    .B1(net35),
    .Y(_0161_));
 sky130_fd_sc_hd__nand4_1 _1724_ (.A(_0274_),
    .B(_0277_),
    .C(\state[2] ),
    .D(\state[0] ),
    .Y(_0192_));
 sky130_fd_sc_hd__nor2_1 _1725_ (.A(\count[0] ),
    .B(_0192_),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_1 _1726_ (.A(_0037_),
    .Y(_0193_));
 sky130_fd_sc_hd__nor2_1 _1727_ (.A(_0193_),
    .B(_0192_),
    .Y(_0163_));
 sky130_fd_sc_hd__xnor2_1 _1728_ (.A(_0036_),
    .B(\count[2] ),
    .Y(_0194_));
 sky130_fd_sc_hd__nor2_1 _1729_ (.A(_0194_),
    .B(_0192_),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_1 _1730_ (.A(\IR[28] ),
    .Y(_0195_));
 sky130_fd_sc_hd__a211oi_1 _1731_ (.A1(_0195_),
    .A2(zero),
    .B1(_0275_),
    .C1(\IR[27] ),
    .Y(_0196_));
 sky130_fd_sc_hd__o21ai_0 _1732_ (.A1(_0414_),
    .A2(_0196_),
    .B1(_0274_),
    .Y(_0197_));
 sky130_fd_sc_hd__a21oi_1 _1733_ (.A1(_0179_),
    .A2(_0414_),
    .B1(_0197_),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_1 _1734_ (.A(\state[2] ),
    .Y(_0198_));
 sky130_fd_sc_hd__nand2_1 _1735_ (.A(_0198_),
    .B(_0174_),
    .Y(_0199_));
 sky130_fd_sc_hd__nand2_1 _1736_ (.A(_0277_),
    .B(\state[2] ),
    .Y(_0200_));
 sky130_fd_sc_hd__a21oi_1 _1737_ (.A1(\state[2] ),
    .A2(\state[1] ),
    .B1(net35),
    .Y(_0201_));
 sky130_fd_sc_hd__nand3_1 _1738_ (.A(_0174_),
    .B(\state[2] ),
    .C(stop),
    .Y(_0202_));
 sky130_fd_sc_hd__nand2_1 _1739_ (.A(_0201_),
    .B(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__a21oi_1 _1740_ (.A1(_0199_),
    .A2(_0200_),
    .B1(_0203_),
    .Y(_0166_));
 sky130_fd_sc_hd__nor2_1 _1741_ (.A(\count[2] ),
    .B(_0198_),
    .Y(_0204_));
 sky130_fd_sc_hd__nor3_1 _1742_ (.A(net35),
    .B(_0908_),
    .C(_0204_),
    .Y(_0167_));
 sky130_fd_sc_hd__nand2_1 _1743_ (.A(_0204_),
    .B(\state[0] ),
    .Y(_0205_));
 sky130_fd_sc_hd__nand3_1 _1744_ (.A(_0205_),
    .B(_0277_),
    .C(_0202_),
    .Y(_0206_));
 sky130_fd_sc_hd__nand2_1 _1745_ (.A(_0206_),
    .B(_0201_),
    .Y(_0207_));
 sky130_fd_sc_hd__inv_1 _1746_ (.A(_0207_),
    .Y(_0168_));
 sky130_fd_sc_hd__nand3_1 _1747_ (.A(\IR[30] ),
    .B(\IR[27] ),
    .C(\IR[28] ),
    .Y(_0208_));
 sky130_fd_sc_hd__o21ai_0 _1748_ (.A1(stop),
    .A2(_0278_),
    .B1(_0274_),
    .Y(_0209_));
 sky130_fd_sc_hd__a21oi_1 _1749_ (.A1(_0278_),
    .A2(_0208_),
    .B1(_0209_),
    .Y(_0169_));
 sky130_fd_sc_hd__nand2_1 _1750_ (.A(_0904_),
    .B(_0905_),
    .Y(_0210_));
 sky130_fd_sc_hd__nand2_1 _1751_ (.A(_0832_),
    .B(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand3_1 _1752_ (.A(_0680_),
    .B(_0624_),
    .C(_0681_),
    .Y(_0212_));
 sky130_fd_sc_hd__nand3_1 _1753_ (.A(_0285_),
    .B(_0035_),
    .C(_0043_),
    .Y(_0213_));
 sky130_fd_sc_hd__nor3_1 _1754_ (.A(_0409_),
    .B(_0213_),
    .C(_0446_),
    .Y(_0214_));
 sky130_fd_sc_hd__nand3_1 _1755_ (.A(_0451_),
    .B(_0489_),
    .C(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__nor2_1 _1756_ (.A(_0215_),
    .B(_0545_),
    .Y(_0216_));
 sky130_fd_sc_hd__nand3_1 _1757_ (.A(_0216_),
    .B(_0558_),
    .C(_0583_),
    .Y(_0217_));
 sky130_fd_sc_hd__nor2_1 _1758_ (.A(_0212_),
    .B(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__nor2_1 _1759_ (.A(_0791_),
    .B(_0806_),
    .Y(_0219_));
 sky130_fd_sc_hd__nor2_1 _1760_ (.A(_0725_),
    .B(_0757_),
    .Y(_0220_));
 sky130_fd_sc_hd__nand3_1 _1761_ (.A(_0218_),
    .B(_0219_),
    .C(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__nor2_1 _1762_ (.A(_0211_),
    .B(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__nand2_1 _1763_ (.A(_0849_),
    .B(_0851_),
    .Y(_0223_));
 sky130_fd_sc_hd__nand2_1 _1764_ (.A(_0712_),
    .B(_0714_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _1765_ (.A(_0798_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__nor2_1 _1766_ (.A(_0223_),
    .B(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__nand2_1 _1767_ (.A(_0747_),
    .B(_0748_),
    .Y(_0227_));
 sky130_fd_sc_hd__nand2_1 _1768_ (.A(_0773_),
    .B(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__nor2_1 _1769_ (.A(_0895_),
    .B(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__nand3_1 _1770_ (.A(_0662_),
    .B(_0597_),
    .C(_0551_),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _1771_ (.A(\IR[16] ),
    .B(_0042_),
    .Y(_0231_));
 sky130_fd_sc_hd__nor2_1 _1772_ (.A(_0231_),
    .B(_0409_),
    .Y(_0232_));
 sky130_fd_sc_hd__nand2_1 _1773_ (.A(_0442_),
    .B(_0444_),
    .Y(_0233_));
 sky130_fd_sc_hd__nand3_1 _1774_ (.A(_0232_),
    .B(_0032_),
    .C(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__nor2_1 _1775_ (.A(_0234_),
    .B(_0465_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand2_1 _1776_ (.A(_0512_),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__nor2_1 _1777_ (.A(_0535_),
    .B(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__nand2_1 _1778_ (.A(_0237_),
    .B(_0616_),
    .Y(_0238_));
 sky130_fd_sc_hd__nor2_1 _1779_ (.A(_0230_),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__nand3_1 _1780_ (.A(_0226_),
    .B(_0229_),
    .C(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__nor2_1 _1781_ (.A(_0418_),
    .B(_0414_),
    .Y(_0241_));
 sky130_fd_sc_hd__nand2_1 _1782_ (.A(_0240_),
    .B(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__nor2_1 _1783_ (.A(_0222_),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__nand3_1 _1784_ (.A(_0741_),
    .B(_0670_),
    .C(_0702_),
    .Y(_0244_));
 sky130_fd_sc_hd__nor2_1 _1785_ (.A(_0604_),
    .B(_0629_),
    .Y(_0245_));
 sky130_fd_sc_hd__nand3b_1 _1786_ (.A_N(_0023_),
    .B(\IR[16] ),
    .C(_0039_),
    .Y(_0246_));
 sky130_fd_sc_hd__nor2_1 _1787_ (.A(_0246_),
    .B(_0435_),
    .Y(_0247_));
 sky130_fd_sc_hd__nand3_1 _1788_ (.A(_0479_),
    .B(_0475_),
    .C(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__nor2_1 _1789_ (.A(_0500_),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__nand2_1 _1790_ (.A(_0249_),
    .B(_0531_),
    .Y(_0250_));
 sky130_fd_sc_hd__nor2_1 _1791_ (.A(_0572_),
    .B(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__nand3_1 _1792_ (.A(_0782_),
    .B(_0245_),
    .C(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__nor2_1 _1793_ (.A(_0244_),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__nand2_1 _1794_ (.A(_0823_),
    .B(_0858_),
    .Y(_0254_));
 sky130_fd_sc_hd__nor2_1 _1795_ (.A(_0874_),
    .B(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__nand2_1 _1796_ (.A(_0253_),
    .B(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__nand2_1 _1797_ (.A(_0845_),
    .B(_0886_),
    .Y(_0257_));
 sky130_fd_sc_hd__nand2_1 _1798_ (.A(_0766_),
    .B(_0817_),
    .Y(_0258_));
 sky130_fd_sc_hd__nor2_1 _1799_ (.A(_0257_),
    .B(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__nor2_1 _1800_ (.A(_0564_),
    .B(_0592_),
    .Y(_0260_));
 sky130_fd_sc_hd__nor4_1 _1801_ (.A(\IR[16] ),
    .B(_0417_),
    .C(_0028_),
    .D(_0439_),
    .Y(_0261_));
 sky130_fd_sc_hd__nand3_1 _1802_ (.A(_0261_),
    .B(_0470_),
    .C(_0506_),
    .Y(_0262_));
 sky130_fd_sc_hd__nor2_1 _1803_ (.A(_0523_),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand3_1 _1804_ (.A(_0260_),
    .B(_0639_),
    .C(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__nand2_1 _1805_ (.A(_0735_),
    .B(_0733_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand3_1 _1806_ (.A(_0691_),
    .B(_0265_),
    .C(_0651_),
    .Y(_0266_));
 sky130_fd_sc_hd__nor2_1 _1807_ (.A(_0264_),
    .B(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__nand2_1 _1808_ (.A(_0259_),
    .B(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__nand2_1 _1809_ (.A(_0256_),
    .B(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__nand2_1 _1810_ (.A(_0269_),
    .B(_0409_),
    .Y(_0270_));
 sky130_fd_sc_hd__o21ai_0 _1811_ (.A1(zero),
    .A2(_0241_),
    .B1(_0274_),
    .Y(_0271_));
 sky130_fd_sc_hd__a21oi_1 _1812_ (.A1(_0243_),
    .A2(_0270_),
    .B1(_0271_),
    .Y(_0170_));
 sky130_fd_sc_hd__fa_1 _1813_ (.A(\IR[1] ),
    .B(net47),
    .CIN(_0021_),
    .COUT(_0022_),
    .SUM(_0023_));
 sky130_fd_sc_hd__fa_1 _1814_ (.A(\GPR[0][1] ),
    .B(net47),
    .CIN(_0026_),
    .COUT(_0027_),
    .SUM(_0028_));
 sky130_fd_sc_hd__fa_1 _1815_ (.A(\IR[1] ),
    .B(_0024_),
    .CIN(_0030_),
    .COUT(_0031_),
    .SUM(_0032_));
 sky130_fd_sc_hd__fa_1 _1816_ (.A(\GPR[0][1] ),
    .B(_0024_),
    .CIN(_0033_),
    .COUT(_0034_),
    .SUM(_0035_));
 sky130_fd_sc_hd__ha_1 _1817_ (.A(\count[0] ),
    .B(\count[1] ),
    .COUT(_0036_),
    .SUM(_0037_));
 sky130_fd_sc_hd__ha_1 _1818_ (.A(_0038_),
    .B(\IR[0] ),
    .COUT(_0030_),
    .SUM(_0039_));
 sky130_fd_sc_hd__ha_1 _1819_ (.A(_0040_),
    .B(\IR[0] ),
    .COUT(_0021_),
    .SUM(_0945_));
 sky130_fd_sc_hd__ha_1 _1820_ (.A(_0038_),
    .B(\GPR[0][0] ),
    .COUT(_0033_),
    .SUM(_0041_));
 sky130_fd_sc_hd__ha_1 _1821_ (.A(_0040_),
    .B(\GPR[0][0] ),
    .COUT(_0026_),
    .SUM(_0946_));
 sky130_fd_sc_hd__ha_1 _1822_ (.A(\IR[0] ),
    .B(_0038_),
    .COUT(_0947_),
    .SUM(_0042_));
 sky130_fd_sc_hd__ha_1 _1823_ (.A(\GPR[0][0] ),
    .B(_0038_),
    .COUT(_0948_),
    .SUM(_0043_));
 sky130_fd_sc_hd__ha_1 _1824_ (.A(net47),
    .B(\IR[1] ),
    .COUT(_0044_),
    .SUM(_0045_));
 sky130_fd_sc_hd__ha_1 _1825_ (.A(net47),
    .B(\GPR[0][1] ),
    .COUT(_0046_),
    .SUM(_0047_));
 sky130_fd_sc_hd__ha_1 _1826_ (.A(_0025_),
    .B(net47),
    .COUT(_0048_),
    .SUM(_0049_));
 sky130_fd_sc_hd__ha_1 _1827_ (.A(_0029_),
    .B(net47),
    .COUT(_0050_),
    .SUM(_0051_));
 sky130_fd_sc_hd__ha_1 _1828_ (.A(\GPR[0][2] ),
    .B(_0052_),
    .COUT(_0053_),
    .SUM(_0054_));
 sky130_fd_sc_hd__ha_1 _1829_ (.A(_0055_),
    .B(_0052_),
    .COUT(_0056_),
    .SUM(_0057_));
 sky130_fd_sc_hd__ha_1 _1830_ (.A(\IR[2] ),
    .B(_0052_),
    .COUT(_0058_),
    .SUM(_0949_));
 sky130_fd_sc_hd__ha_1 _1831_ (.A(_0059_),
    .B(_0052_),
    .COUT(_0060_),
    .SUM(_0061_));
 sky130_fd_sc_hd__ha_1 _1832_ (.A(_0062_),
    .B(\GPR[0][3] ),
    .COUT(_0063_),
    .SUM(_0064_));
 sky130_fd_sc_hd__ha_1 _1833_ (.A(_0065_),
    .B(_0062_),
    .COUT(_0066_),
    .SUM(_0067_));
 sky130_fd_sc_hd__ha_1 _1834_ (.A(_0068_),
    .B(\GPR[0][4] ),
    .COUT(_0069_),
    .SUM(_0070_));
 sky130_fd_sc_hd__ha_1 _1835_ (.A(_0071_),
    .B(_0068_),
    .COUT(_0072_),
    .SUM(_0073_));
 sky130_fd_sc_hd__ha_1 _1836_ (.A(\GPR[0][5] ),
    .B(_0074_),
    .COUT(_0075_),
    .SUM(_0076_));
 sky130_fd_sc_hd__ha_1 _1837_ (.A(_0077_),
    .B(_0074_),
    .COUT(_0078_),
    .SUM(_0079_));
 sky130_fd_sc_hd__ha_1 _1838_ (.A(\GPR[0][6] ),
    .B(_0080_),
    .COUT(_0081_),
    .SUM(_0082_));
 sky130_fd_sc_hd__ha_1 _1839_ (.A(_0083_),
    .B(_0080_),
    .COUT(_0084_),
    .SUM(_0085_));
 sky130_fd_sc_hd__ha_1 _1840_ (.A(_0086_),
    .B(\GPR[0][7] ),
    .COUT(_0087_),
    .SUM(_0088_));
 sky130_fd_sc_hd__ha_1 _1841_ (.A(_0086_),
    .B(_0089_),
    .COUT(_0090_),
    .SUM(_0091_));
 sky130_fd_sc_hd__ha_1 _1842_ (.A(_0092_),
    .B(\GPR[0][8] ),
    .COUT(_0093_),
    .SUM(_0094_));
 sky130_fd_sc_hd__ha_1 _1843_ (.A(_0095_),
    .B(_0092_),
    .COUT(_0096_),
    .SUM(_0097_));
 sky130_fd_sc_hd__ha_1 _1844_ (.A(_0098_),
    .B(\GPR[0][9] ),
    .COUT(_0099_),
    .SUM(_0100_));
 sky130_fd_sc_hd__ha_1 _1845_ (.A(_0101_),
    .B(_0098_),
    .COUT(_0102_),
    .SUM(_0103_));
 sky130_fd_sc_hd__ha_1 _1846_ (.A(_0104_),
    .B(\GPR[0][10] ),
    .COUT(_0105_),
    .SUM(_0106_));
 sky130_fd_sc_hd__ha_1 _1847_ (.A(_0107_),
    .B(_0104_),
    .COUT(_0108_),
    .SUM(_0109_));
 sky130_fd_sc_hd__ha_1 _1848_ (.A(_0110_),
    .B(\GPR[0][11] ),
    .COUT(_0111_),
    .SUM(_0112_));
 sky130_fd_sc_hd__ha_1 _1849_ (.A(_0110_),
    .B(_0113_),
    .COUT(_0114_),
    .SUM(_0115_));
 sky130_fd_sc_hd__ha_1 _1850_ (.A(_0116_),
    .B(\GPR[0][12] ),
    .COUT(_0117_),
    .SUM(_0118_));
 sky130_fd_sc_hd__ha_1 _1851_ (.A(_0119_),
    .B(_0116_),
    .COUT(_0120_),
    .SUM(_0121_));
 sky130_fd_sc_hd__ha_1 _1852_ (.A(_0122_),
    .B(\GPR[0][13] ),
    .COUT(_0123_),
    .SUM(_0124_));
 sky130_fd_sc_hd__ha_1 _1853_ (.A(_0125_),
    .B(_0122_),
    .COUT(_0126_),
    .SUM(_0127_));
 sky130_fd_sc_hd__ha_1 _1854_ (.A(_0128_),
    .B(_0129_),
    .COUT(_0130_),
    .SUM(_0131_));
 sky130_fd_sc_hd__ha_1 _1855_ (.A(_0129_),
    .B(_0128_),
    .COUT(_0950_),
    .SUM(_0132_));
 sky130_fd_sc_hd__ha_1 _1856_ (.A(\GPR[0][14] ),
    .B(_0128_),
    .COUT(_0133_),
    .SUM(_0951_));
 sky130_fd_sc_hd__ha_1 _1857_ (.A(_0134_),
    .B(_0135_),
    .COUT(_0136_),
    .SUM(_0137_));
 sky130_fd_sc_hd__ha_1 _1858_ (.A(_0134_),
    .B(\PC[1] ),
    .COUT(_0138_),
    .SUM(_0952_));
 sky130_fd_sc_hd__ha_1 _1859_ (.A(_0134_),
    .B(\PC[1] ),
    .COUT(_0139_),
    .SUM(_0953_));
 sky130_fd_sc_hd__ha_1 _1860_ (.A(\PC[0] ),
    .B(_0135_),
    .COUT(_0140_),
    .SUM(_0954_));
 sky130_fd_sc_hd__ha_1 _1861_ (.A(\PC[0] ),
    .B(\PC[1] ),
    .COUT(_0955_),
    .SUM(_0956_));
 sky130_fd_sc_hd__ha_1 _1862_ (.A(\PC[2] ),
    .B(_0955_),
    .COUT(_0141_),
    .SUM(_0142_));
 sky130_fd_sc_hd__ha_1 _1863_ (.A(_0135_),
    .B(\PC[2] ),
    .COUT(_0143_),
    .SUM(_0144_));
 sky130_fd_sc_hd__ha_1 _1864_ (.A(\PC[1] ),
    .B(\PC[2] ),
    .COUT(_0145_),
    .SUM(_0957_));
 sky130_fd_sc_hd__inv_6 clkload6 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload5 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload4 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__buf_4 place49 (.A(\IR[18] ),
    .X(net48));
 sky130_fd_sc_hd__buf_4 place48 (.A(_0020_),
    .X(net47));
 sky130_fd_sc_hd__buf_4 place43 (.A(_0016_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_4 place50 (.A(\IR[17] ),
    .X(net49));
 sky130_fd_sc_hd__buf_4 place47 (.A(_0415_),
    .X(net46));
 sky130_fd_sc_hd__buf_4 place46 (.A(_0019_),
    .X(net45));
 sky130_fd_sc_hd__buf_4 place45 (.A(_0018_),
    .X(net44));
 sky130_fd_sc_hd__buf_4 place44 (.A(_0017_),
    .X(net43));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input36 (.A(sys_rst),
    .X(net35));
 sky130_fd_sc_hd__dfxtp_1 \count[0]$_SDFF_PP0_  (.D(_0162_),
    .Q(\count[0] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \count[1]$_SDFF_PP0_  (.D(_0163_),
    .Q(\count[1] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \count[2]$_SDFF_PP0_  (.D(_0164_),
    .Q(\count[2] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \jmp_flag$_SDFFE_PP0P_  (.D(_0165_),
    .Q(jmp_flag),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \state[0]$_SDFF_PP0_  (.D(_0166_),
    .Q(\state[0] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \state[1]$_SDFF_PP0_  (.D(_0167_),
    .Q(\state[1] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \state[2]$_SDFF_PP0_  (.D(_0168_),
    .Q(\state[2] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \stop$_SDFFE_PP0P_  (.D(_0169_),
    .Q(stop),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \zero$_SDFFE_PP0P_  (.D(_0170_),
    .Q(zero),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__conb_1 _1866__1 (.LO(net));
 sky130_fd_sc_hd__conb_1 _1867__2 (.LO(net1));
 sky130_fd_sc_hd__conb_1 _1868__3 (.LO(net2));
 sky130_fd_sc_hd__conb_1 _1869__4 (.LO(net3));
 sky130_fd_sc_hd__conb_1 _1870__5 (.LO(net4));
 sky130_fd_sc_hd__conb_1 _1871__6 (.LO(net5));
 sky130_fd_sc_hd__conb_1 _1872__7 (.LO(net6));
 sky130_fd_sc_hd__conb_1 _1873__8 (.LO(net7));
 sky130_fd_sc_hd__conb_1 _1874__9 (.LO(net8));
 sky130_fd_sc_hd__conb_1 _1875__10 (.LO(net9));
 sky130_fd_sc_hd__conb_1 _1876__11 (.LO(net10));
 sky130_fd_sc_hd__conb_1 _1877__12 (.LO(net11));
 sky130_fd_sc_hd__conb_1 _1878__13 (.LO(net12));
 sky130_fd_sc_hd__conb_1 _1879__14 (.LO(net13));
 sky130_fd_sc_hd__conb_1 _1880__15 (.LO(net14));
 sky130_fd_sc_hd__conb_1 _1881__16 (.LO(net15));
 sky130_fd_sc_hd__conb_1 _1882__17 (.LO(net16));
 sky130_fd_sc_hd__conb_1 _1883__18 (.LO(net17));
 sky130_fd_sc_hd__conb_1 _1884__19 (.LO(net18));
 sky130_fd_sc_hd__conb_1 _1885__20 (.LO(dout[0]));
 sky130_fd_sc_hd__conb_1 _1886__21 (.LO(dout[1]));
 sky130_fd_sc_hd__conb_1 _1887__22 (.LO(dout[2]));
 sky130_fd_sc_hd__conb_1 _1888__23 (.LO(dout[3]));
 sky130_fd_sc_hd__conb_1 _1889__24 (.LO(dout[4]));
 sky130_fd_sc_hd__conb_1 _1890__25 (.LO(dout[5]));
 sky130_fd_sc_hd__conb_1 _1891__26 (.LO(dout[6]));
 sky130_fd_sc_hd__conb_1 _1892__27 (.LO(dout[7]));
 sky130_fd_sc_hd__conb_1 _1893__28 (.LO(dout[8]));
 sky130_fd_sc_hd__conb_1 _1894__29 (.LO(dout[9]));
 sky130_fd_sc_hd__conb_1 _1895__30 (.LO(dout[10]));
 sky130_fd_sc_hd__conb_1 _1896__31 (.LO(dout[11]));
 sky130_fd_sc_hd__conb_1 _1897__32 (.LO(dout[12]));
 sky130_fd_sc_hd__conb_1 _1898__33 (.LO(dout[13]));
 sky130_fd_sc_hd__conb_1 _1899__34 (.LO(dout[14]));
 sky130_fd_sc_hd__conb_1 _1900__35 (.LO(dout[15]));
endmodule
